.title <test_1R_cb_4x4_2f>


** Includes **


** Load models **
.hdl ../models/rram_wp.va

** Options **
.option post=2

** Parameters **


** Probes **


** Sub-circuits **
.subckt CELL r1 r2 c1 c2 gap
Ccell r1 c1 1f
Rr r1 r2 0.18
Cr r2 gnd 1.08e-13
Rc c1 c2 0.18
Cc c2 gnd 1.08e-13
X1 r1 c1 gap RRAM_v0 
.ends CELL


** Crossbar instantiation **
Xcell_0_0 row_0_0 row_0_1 col_0_0 col_1_0 gap_0_0 CELL
.nodeset gap_0_0 0.85
Xcell_0_1 row_0_1 row_0_2 col_0_1 col_1_1 gap_0_1 CELL
.nodeset gap_0_1 0.85
Xcell_0_2 row_0_2 row_0_3 col_0_2 col_1_2 gap_0_2 CELL
.nodeset gap_0_2 0.85
Xcell_0_3 row_0_3 row_0_4 col_0_3 col_1_3 gap_0_3 CELL
.nodeset gap_0_3 0.85
Xcell_1_0 row_1_0 row_1_1 col_1_0 col_2_0 gap_1_0 CELL
.nodeset gap_1_0 0.85
Xcell_1_1 row_1_1 row_1_2 col_1_1 col_2_1 gap_1_1 CELL
.nodeset gap_1_1 0.85
Xcell_1_2 row_1_2 row_1_3 col_1_2 col_2_2 gap_1_2 CELL
.nodeset gap_1_2 0.85
Xcell_1_3 row_1_3 row_1_4 col_1_3 col_2_3 gap_1_3 CELL
.nodeset gap_1_3 0.85
Xcell_2_0 row_2_0 row_2_1 col_2_0 col_3_0 gap_2_0 CELL
.nodeset gap_2_0 0.85
Xcell_2_1 row_2_1 row_2_2 col_2_1 col_3_1 gap_2_1 CELL
.nodeset gap_2_1 0.85
Xcell_2_2 row_2_2 row_2_3 col_2_2 col_3_2 gap_2_2 CELL
.nodeset gap_2_2 0.85
Xcell_2_3 row_2_3 row_2_4 col_2_3 col_3_3 gap_2_3 CELL
.nodeset gap_2_3 0.85
Xcell_3_0 row_3_0 row_3_1 col_3_0 col_4_0 gap_3_0 CELL
.nodeset gap_3_0 0.85
Xcell_3_1 row_3_1 row_3_2 col_3_1 col_4_1 gap_3_1 CELL
.nodeset gap_3_1 0.85
Xcell_3_2 row_3_2 row_3_3 col_3_2 col_4_2 gap_3_2 CELL
.nodeset gap_3_2 0.85
Xcell_3_3 row_3_3 row_3_4 col_3_3 col_4_3 gap_3_3 CELL
.nodeset gap_3_3 0.85


** PWL voltage waveforms **
Vrow_0 row_0_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 0.2            4.9e-06 0.2          5e-06 0              5.9e-06 0            6e-06 0.2            6.9e-06 0.2          7e-06 0              7.9e-06 0            8e-06 0.2            8.9e-06 0.2          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 0            3.69e-05 0           3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 0              4.09e-05 0           4.1e-05 0            4.19e-05 0           4.2e-05 0.75         4.29e-05 0.75        4.3e-05 0            4.39e-05 0           4.4e-05 0.75         4.49e-05 0.75        4.5e-05 0            4.59e-05 0           4.6e-05 0.75         4.69e-05 0.75        4.7e-05 0            4.79e-05 0           4.8e-05 0.75         4.89e-05 0.75        4.9e-05 0            4.99e-05 0           5e-05 0.75           5.09e-05 0.75        5.1e-05 0            5.19e-05 0           5.2e-05 0.75         5.29e-05 0.75        5.3e-05 0            5.39e-05 0           5.4e-05 0.75         5.49e-05 0.75        5.5e-05 0            5.59e-05 0           5.6e-05 0.75         5.69e-05 0.75        5.7e-05 0            5.79e-05 0           5.8e-05 0.75         5.89e-05 0.75        5.9e-05 0            5.99e-05 0           6e-05 0.75           6.09e-05 0.75        6.1e-05 0            6.19e-05 0           6.2e-05 0.75         6.29e-05 0.75        6.3e-05 0            6.39e-05 0           6.4e-05 0.75         6.49e-05 0.75        6.5e-05 0            6.59e-05 0           6.6e-05 0.2          6.69e-05 0.2         6.7e-05 0            6.79e-05 0           6.8e-05 0.2          6.89e-05 0.2         6.9e-05 0            6.99e-05 0           7e-05 0.2            7.09e-05 0.2         7.1e-05 0            7.19e-05 0           7.2e-05 0.2          7.29e-05 0.2         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0            9.89e-05 0           9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 0           0.0001029 0          0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 0.75        0.0001069 0.75       0.000107 0           0.0001079 0          0.000108 0.75        0.0001089 0.75       0.000109 0           0.0001099 0          0.00011 0.75         0.0001109 0.75       0.000111 0           0.0001119 0          0.000112 0.75        0.0001129 0.75       0.000113 0           0.0001139 0          0.000114 0.75        0.0001149 0.75       0.000115 0           0.0001159 0          0.000116 0.75        0.0001169 0.75       0.000117 0           0.0001179 0          0.000118 0.75        0.0001189 0.75       0.000119 0           0.0001199 0          0.00012 0.75         0.0001209 0.75       0.000121 0           0.0001219 0          0.000122 0.75        0.0001229 0.75       0.000123 0           0.0001239 0          0.000124 0.75        0.0001249 0.75       0.000125 0           0.0001259 0          0.000126 0.75        0.0001269 0.75       0.000127 0           0.0001279 0          0.000128 0.75        0.0001289 0.75       0.000129 0           0.0001299 0          0.00013 0.2          0.0001309 0.2        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 0.2         0.0001349 0.2        0.000135 0           0.0001359 0          0.000136 0.2         0.0001369 0.2        0.000137 0           0.0001379 0          0.000138 0.1         0.0001389 0.1        0.000139 0           0.0001399 0          0.00014 0.1          0.0001409 0.1        0.000141 0           0.0001419 0          0.000142 0.1         0.0001429 0.1        0.000143 0           0.0001439 0          0.000144 0.1         0.0001449 0.1        0.000145 0           0.0001459 0          0.000146 0.1         0.0001469 0.1        0.000147 0           0.0001479 0          0.000148 0.1         0.0001489 0.1        0.000149 0           0.0001499 0          0.00015 0.1          0.0001509 0.1        0.000151 0           0.0001519 0          0.000152 0.1         0.0001529 0.1        0.000153 0           0.0001539 0          0.000154 0.1         0.0001549 0.1        0.000155 0           0.0001559 0          0.000156 0.1         0.0001569 0.1        0.000157 0           0.0001579 0          0.000158 0.1         0.0001589 0.1        0.000159 0           0.0001599 0          0.00016 0.1          0.0001609 0.1        0.000161 0           0.0001619 0         )
Vrow_1 row_1_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.2            1.09e-05 0.2         1.1e-05 0            1.19e-05 0           1.2e-05 0.2          1.29e-05 0.2         1.3e-05 0            1.39e-05 0           1.4e-05 0.2          1.49e-05 0.2         1.5e-05 0            1.59e-05 0           1.6e-05 0.2          1.69e-05 0.2         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.75         3.49e-05 0.75        3.5e-05 0            3.59e-05 0           3.6e-05 0.75         3.69e-05 0.75        3.7e-05 0            3.79e-05 0           3.8e-05 0.75         3.89e-05 0.75        3.9e-05 0            3.99e-05 0           4e-05 0.75           4.09e-05 0.75        4.1e-05 0            4.19e-05 0           4.2e-05 0            4.29e-05 0           4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 0            4.69e-05 0           4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 0.75           5.09e-05 0.75        5.1e-05 0            5.19e-05 0           5.2e-05 0.75         5.29e-05 0.75        5.3e-05 0            5.39e-05 0           5.4e-05 0.75         5.49e-05 0.75        5.5e-05 0            5.59e-05 0           5.6e-05 0.75         5.69e-05 0.75        5.7e-05 0            5.79e-05 0           5.8e-05 0.75         5.89e-05 0.75        5.9e-05 0            5.99e-05 0           6e-05 0.75           6.09e-05 0.75        6.1e-05 0            6.19e-05 0           6.2e-05 0.75         6.29e-05 0.75        6.3e-05 0            6.39e-05 0           6.4e-05 0.75         6.49e-05 0.75        6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.2          7.49e-05 0.2         7.5e-05 0            7.59e-05 0           7.6e-05 0.2          7.69e-05 0.2         7.7e-05 0            7.79e-05 0           7.8e-05 0.2          7.89e-05 0.2         7.9e-05 0            7.99e-05 0           8e-05 0.2            8.09e-05 0.2         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.75         9.89e-05 0.75        9.9e-05 0            9.99e-05 0           0.0001 0.75          0.0001009 0.75       0.000101 0           0.0001019 0          0.000102 0.75        0.0001029 0.75       0.000103 0           0.0001039 0          0.000104 0.75        0.0001049 0.75       0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 0           0.0001089 0          0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 0           0.0001129 0          0.000113 0           0.0001139 0          0.000114 0.75        0.0001149 0.75       0.000115 0           0.0001159 0          0.000116 0.75        0.0001169 0.75       0.000117 0           0.0001179 0          0.000118 0.75        0.0001189 0.75       0.000119 0           0.0001199 0          0.00012 0.75         0.0001209 0.75       0.000121 0           0.0001219 0          0.000122 0.75        0.0001229 0.75       0.000123 0           0.0001239 0          0.000124 0.75        0.0001249 0.75       0.000125 0           0.0001259 0          0.000126 0.75        0.0001269 0.75       0.000127 0           0.0001279 0          0.000128 0.75        0.0001289 0.75       0.000129 0           0.0001299 0          0.00013 0.1          0.0001309 0.1        0.000131 0           0.0001319 0          0.000132 0.1         0.0001329 0.1        0.000133 0           0.0001339 0          0.000134 0.1         0.0001349 0.1        0.000135 0           0.0001359 0          0.000136 0.1         0.0001369 0.1        0.000137 0           0.0001379 0          0.000138 0.2         0.0001389 0.2        0.000139 0           0.0001399 0          0.00014 0.2          0.0001409 0.2        0.000141 0           0.0001419 0          0.000142 0.2         0.0001429 0.2        0.000143 0           0.0001439 0          0.000144 0.2         0.0001449 0.2        0.000145 0           0.0001459 0          0.000146 0.1         0.0001469 0.1        0.000147 0           0.0001479 0          0.000148 0.1         0.0001489 0.1        0.000149 0           0.0001499 0          0.00015 0.1          0.0001509 0.1        0.000151 0           0.0001519 0          0.000152 0.1         0.0001529 0.1        0.000153 0           0.0001539 0          0.000154 0.1         0.0001549 0.1        0.000155 0           0.0001559 0          0.000156 0.1         0.0001569 0.1        0.000157 0           0.0001579 0          0.000158 0.1         0.0001589 0.1        0.000159 0           0.0001599 0          0.00016 0.1          0.0001609 0.1        0.000161 0           0.0001619 0         )
Vrow_2 row_2_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.2          1.89e-05 0.2         1.9e-05 0            1.99e-05 0           2e-05 0.2            2.09e-05 0.2         2.1e-05 0            2.19e-05 0           2.2e-05 0.2          2.29e-05 0.2         2.3e-05 0            2.39e-05 0           2.4e-05 0.2          2.49e-05 0.2         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.75         3.49e-05 0.75        3.5e-05 0            3.59e-05 0           3.6e-05 0.75         3.69e-05 0.75        3.7e-05 0            3.79e-05 0           3.8e-05 0.75         3.89e-05 0.75        3.9e-05 0            3.99e-05 0           4e-05 0.75           4.09e-05 0.75        4.1e-05 0            4.19e-05 0           4.2e-05 0.75         4.29e-05 0.75        4.3e-05 0            4.39e-05 0           4.4e-05 0.75         4.49e-05 0.75        4.5e-05 0            4.59e-05 0           4.6e-05 0.75         4.69e-05 0.75        4.7e-05 0            4.79e-05 0           4.8e-05 0.75         4.89e-05 0.75        4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 0            5.29e-05 0           5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 0            5.69e-05 0           5.7e-05 0            5.79e-05 0           5.8e-05 0.75         5.89e-05 0.75        5.9e-05 0            5.99e-05 0           6e-05 0.75           6.09e-05 0.75        6.1e-05 0            6.19e-05 0           6.2e-05 0.75         6.29e-05 0.75        6.3e-05 0            6.39e-05 0           6.4e-05 0.75         6.49e-05 0.75        6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.2          8.29e-05 0.2         8.3e-05 0            8.39e-05 0           8.4e-05 0.2          8.49e-05 0.2         8.5e-05 0            8.59e-05 0           8.6e-05 0.2          8.69e-05 0.2         8.7e-05 0            8.79e-05 0           8.8e-05 0.2          8.89e-05 0.2         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.75         9.89e-05 0.75        9.9e-05 0            9.99e-05 0           0.0001 0.75          0.0001009 0.75       0.000101 0           0.0001019 0          0.000102 0.75        0.0001029 0.75       0.000103 0           0.0001039 0          0.000104 0.75        0.0001049 0.75       0.000105 0           0.0001059 0          0.000106 0.75        0.0001069 0.75       0.000107 0           0.0001079 0          0.000108 0.75        0.0001089 0.75       0.000109 0           0.0001099 0          0.00011 0.75         0.0001109 0.75       0.000111 0           0.0001119 0          0.000112 0.75        0.0001129 0.75       0.000113 0           0.0001139 0          0.000114 0           0.0001149 0          0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 0           0.0001189 0          0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 0.75        0.0001229 0.75       0.000123 0           0.0001239 0          0.000124 0.75        0.0001249 0.75       0.000125 0           0.0001259 0          0.000126 0.75        0.0001269 0.75       0.000127 0           0.0001279 0          0.000128 0.75        0.0001289 0.75       0.000129 0           0.0001299 0          0.00013 0.1          0.0001309 0.1        0.000131 0           0.0001319 0          0.000132 0.1         0.0001329 0.1        0.000133 0           0.0001339 0          0.000134 0.1         0.0001349 0.1        0.000135 0           0.0001359 0          0.000136 0.1         0.0001369 0.1        0.000137 0           0.0001379 0          0.000138 0.1         0.0001389 0.1        0.000139 0           0.0001399 0          0.00014 0.1          0.0001409 0.1        0.000141 0           0.0001419 0          0.000142 0.1         0.0001429 0.1        0.000143 0           0.0001439 0          0.000144 0.1         0.0001449 0.1        0.000145 0           0.0001459 0          0.000146 0.2         0.0001469 0.2        0.000147 0           0.0001479 0          0.000148 0.2         0.0001489 0.2        0.000149 0           0.0001499 0          0.00015 0.2          0.0001509 0.2        0.000151 0           0.0001519 0          0.000152 0.2         0.0001529 0.2        0.000153 0           0.0001539 0          0.000154 0.1         0.0001549 0.1        0.000155 0           0.0001559 0          0.000156 0.1         0.0001569 0.1        0.000157 0           0.0001579 0          0.000158 0.1         0.0001589 0.1        0.000159 0           0.0001599 0          0.00016 0.1          0.0001609 0.1        0.000161 0           0.0001619 0         )
Vrow_3 row_3_0 0 PWLZ(0 0                  9e-07 0              1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.2          2.69e-05 0.2         2.7e-05 0            2.79e-05 0           2.8e-05 0.2          2.89e-05 0.2         2.9e-05 0            2.99e-05 0           3e-05 0.2            3.09e-05 0.2         3.1e-05 0            3.19e-05 0           3.2e-05 0.2          3.29e-05 0.2         3.3e-05 0            3.39e-05 0           3.4e-05 0.75         3.49e-05 0.75        3.5e-05 0            3.59e-05 0           3.6e-05 0.75         3.69e-05 0.75        3.7e-05 0            3.79e-05 0           3.8e-05 0.75         3.89e-05 0.75        3.9e-05 0            3.99e-05 0           4e-05 0.75           4.09e-05 0.75        4.1e-05 0            4.19e-05 0           4.2e-05 0.75         4.29e-05 0.75        4.3e-05 0            4.39e-05 0           4.4e-05 0.75         4.49e-05 0.75        4.5e-05 0            4.59e-05 0           4.6e-05 0.75         4.69e-05 0.75        4.7e-05 0            4.79e-05 0           4.8e-05 0.75         4.89e-05 0.75        4.9e-05 0            4.99e-05 0           5e-05 0.75           5.09e-05 0.75        5.1e-05 0            5.19e-05 0           5.2e-05 0.75         5.29e-05 0.75        5.3e-05 0            5.39e-05 0           5.4e-05 0.75         5.49e-05 0.75        5.5e-05 0            5.59e-05 0           5.6e-05 0.75         5.69e-05 0.75        5.7e-05 0            5.79e-05 0           5.8e-05 0            5.89e-05 0           5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 0            6.29e-05 0           6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.2            9.09e-05 0.2         9.1e-05 0            9.19e-05 0           9.2e-05 0.2          9.29e-05 0.2         9.3e-05 0            9.39e-05 0           9.4e-05 0.2          9.49e-05 0.2         9.5e-05 0            9.59e-05 0           9.6e-05 0.2          9.69e-05 0.2         9.7e-05 0            9.79e-05 0           9.8e-05 0.75         9.89e-05 0.75        9.9e-05 0            9.99e-05 0           0.0001 0.75          0.0001009 0.75       0.000101 0           0.0001019 0          0.000102 0.75        0.0001029 0.75       0.000103 0           0.0001039 0          0.000104 0.75        0.0001049 0.75       0.000105 0           0.0001059 0          0.000106 0.75        0.0001069 0.75       0.000107 0           0.0001079 0          0.000108 0.75        0.0001089 0.75       0.000109 0           0.0001099 0          0.00011 0.75         0.0001109 0.75       0.000111 0           0.0001119 0          0.000112 0.75        0.0001129 0.75       0.000113 0           0.0001139 0          0.000114 0.75        0.0001149 0.75       0.000115 0           0.0001159 0          0.000116 0.75        0.0001169 0.75       0.000117 0           0.0001179 0          0.000118 0.75        0.0001189 0.75       0.000119 0           0.0001199 0          0.00012 0.75         0.0001209 0.75       0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 0           0.0001249 0          0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 0           0.0001289 0          0.000129 0           0.0001299 0          0.00013 0.1          0.0001309 0.1        0.000131 0           0.0001319 0          0.000132 0.1         0.0001329 0.1        0.000133 0           0.0001339 0          0.000134 0.1         0.0001349 0.1        0.000135 0           0.0001359 0          0.000136 0.1         0.0001369 0.1        0.000137 0           0.0001379 0          0.000138 0.1         0.0001389 0.1        0.000139 0           0.0001399 0          0.00014 0.1          0.0001409 0.1        0.000141 0           0.0001419 0          0.000142 0.1         0.0001429 0.1        0.000143 0           0.0001439 0          0.000144 0.1         0.0001449 0.1        0.000145 0           0.0001459 0          0.000146 0.1         0.0001469 0.1        0.000147 0           0.0001479 0          0.000148 0.1         0.0001489 0.1        0.000149 0           0.0001499 0          0.00015 0.1          0.0001509 0.1        0.000151 0           0.0001519 0          0.000152 0.1         0.0001529 0.1        0.000153 0           0.0001539 0          0.000154 0.2         0.0001549 0.2        0.000155 0           0.0001559 0          0.000156 0.2         0.0001569 0.2        0.000157 0           0.0001579 0          0.000158 0.2         0.0001589 0.2        0.000159 0           0.0001599 0          0.00016 0.2          0.0001609 0.2        0.000161 0           0.0001619 0         )
Vcol_0 col_0_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0              1.09e-05 0           1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0            1.89e-05 0           1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0            2.69e-05 0           2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0            3.49e-05 0           3.5e-05 0            3.59e-05 0           3.6e-05 0.75         3.69e-05 0.75        3.7e-05 0            3.79e-05 0           3.8e-05 0.75         3.89e-05 0.75        3.9e-05 0            3.99e-05 0           4e-05 0.75           4.09e-05 0.75        4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 0.75         4.49e-05 0.75        4.5e-05 0            4.59e-05 0           4.6e-05 0.75         4.69e-05 0.75        4.7e-05 0            4.79e-05 0           4.8e-05 0.75         4.89e-05 0.75        4.9e-05 0            4.99e-05 0           5e-05 0              5.09e-05 0           5.1e-05 0            5.19e-05 0           5.2e-05 0.75         5.29e-05 0.75        5.3e-05 0            5.39e-05 0           5.4e-05 0.75         5.49e-05 0.75        5.5e-05 0            5.59e-05 0           5.6e-05 0.75         5.69e-05 0.75        5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 0.75           6.09e-05 0.75        6.1e-05 0            6.19e-05 0           6.2e-05 0.75         6.29e-05 0.75        6.3e-05 0            6.39e-05 0           6.4e-05 0.75         6.49e-05 0.75        6.5e-05 0            6.59e-05 0           6.6e-05 0            6.69e-05 0           6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0            7.49e-05 0           7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0            8.29e-05 0           8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0              9.09e-05 0           9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 0.75          0.0001009 0.75       0.000101 0           0.0001019 0          0.000102 0.75        0.0001029 0.75       0.000103 0           0.0001039 0          0.000104 0.75        0.0001049 0.75       0.000105 0           0.0001059 0          0.000106 0           0.0001069 0          0.000107 0           0.0001079 0          0.000108 0.75        0.0001089 0.75       0.000109 0           0.0001099 0          0.00011 0.75         0.0001109 0.75       0.000111 0           0.0001119 0          0.000112 0.75        0.0001129 0.75       0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 0.75        0.0001169 0.75       0.000117 0           0.0001179 0          0.000118 0.75        0.0001189 0.75       0.000119 0           0.0001199 0          0.00012 0.75         0.0001209 0.75       0.000121 0           0.0001219 0          0.000122 0           0.0001229 0          0.000123 0           0.0001239 0          0.000124 0.75        0.0001249 0.75       0.000125 0           0.0001259 0          0.000126 0.75        0.0001269 0.75       0.000127 0           0.0001279 0          0.000128 0.75        0.0001289 0.75       0.000129 0           0.0001299 0          0.00013 0            0.0001309 0          0.000131 0           0.0001319 0          0.000132 0.1         0.0001329 0.1        0.000133 0           0.0001339 0          0.000134 0.1         0.0001349 0.1        0.000135 0           0.0001359 0          0.000136 0.1         0.0001369 0.1        0.000137 0           0.0001379 0          0.000138 0           0.0001389 0          0.000139 0           0.0001399 0          0.00014 0.1          0.0001409 0.1        0.000141 0           0.0001419 0          0.000142 0.1         0.0001429 0.1        0.000143 0           0.0001439 0          0.000144 0.1         0.0001449 0.1        0.000145 0           0.0001459 0          0.000146 0           0.0001469 0          0.000147 0           0.0001479 0          0.000148 0.1         0.0001489 0.1        0.000149 0           0.0001499 0          0.00015 0.1          0.0001509 0.1        0.000151 0           0.0001519 0          0.000152 0.1         0.0001529 0.1        0.000153 0           0.0001539 0          0.000154 0           0.0001549 0          0.000155 0           0.0001559 0          0.000156 0.1         0.0001569 0.1        0.000157 0           0.0001579 0          0.000158 0.1         0.0001589 0.1        0.000159 0           0.0001599 0          0.00016 0.1          0.0001609 0.1        0.000161 0           0.0001619 0         )
Vcol_1 col_0_1 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0              4.9e-06 0            5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0            1.29e-05 0           1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0              2.09e-05 0           2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0            2.89e-05 0           2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.75         3.49e-05 0.75        3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 0.75         3.89e-05 0.75        3.9e-05 0            3.99e-05 0           4e-05 0.75           4.09e-05 0.75        4.1e-05 0            4.19e-05 0           4.2e-05 0.75         4.29e-05 0.75        4.3e-05 0            4.39e-05 0           4.4e-05 0            4.49e-05 0           4.5e-05 0            4.59e-05 0           4.6e-05 0.75         4.69e-05 0.75        4.7e-05 0            4.79e-05 0           4.8e-05 0.75         4.89e-05 0.75        4.9e-05 0            4.99e-05 0           5e-05 0.75           5.09e-05 0.75        5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 0.75         5.49e-05 0.75        5.5e-05 0            5.59e-05 0           5.6e-05 0.75         5.69e-05 0.75        5.7e-05 0            5.79e-05 0           5.8e-05 0.75         5.89e-05 0.75        5.9e-05 0            5.99e-05 0           6e-05 0              6.09e-05 0           6.1e-05 0            6.19e-05 0           6.2e-05 0.75         6.29e-05 0.75        6.3e-05 0            6.39e-05 0           6.4e-05 0.75         6.49e-05 0.75        6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0            6.89e-05 0           6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0            7.69e-05 0           7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0            8.49e-05 0           8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0            9.29e-05 0           9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.75         9.89e-05 0.75        9.9e-05 0            9.99e-05 0           0.0001 0             0.0001009 0          0.000101 0           0.0001019 0          0.000102 0.75        0.0001029 0.75       0.000103 0           0.0001039 0          0.000104 0.75        0.0001049 0.75       0.000105 0           0.0001059 0          0.000106 0.75        0.0001069 0.75       0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 0.75         0.0001109 0.75       0.000111 0           0.0001119 0          0.000112 0.75        0.0001129 0.75       0.000113 0           0.0001139 0          0.000114 0.75        0.0001149 0.75       0.000115 0           0.0001159 0          0.000116 0           0.0001169 0          0.000117 0           0.0001179 0          0.000118 0.75        0.0001189 0.75       0.000119 0           0.0001199 0          0.00012 0.75         0.0001209 0.75       0.000121 0           0.0001219 0          0.000122 0.75        0.0001229 0.75       0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 0.75        0.0001269 0.75       0.000127 0           0.0001279 0          0.000128 0.75        0.0001289 0.75       0.000129 0           0.0001299 0          0.00013 0.1          0.0001309 0.1        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 0.1         0.0001349 0.1        0.000135 0           0.0001359 0          0.000136 0.1         0.0001369 0.1        0.000137 0           0.0001379 0          0.000138 0.1         0.0001389 0.1        0.000139 0           0.0001399 0          0.00014 0            0.0001409 0          0.000141 0           0.0001419 0          0.000142 0.1         0.0001429 0.1        0.000143 0           0.0001439 0          0.000144 0.1         0.0001449 0.1        0.000145 0           0.0001459 0          0.000146 0.1         0.0001469 0.1        0.000147 0           0.0001479 0          0.000148 0           0.0001489 0          0.000149 0           0.0001499 0          0.00015 0.1          0.0001509 0.1        0.000151 0           0.0001519 0          0.000152 0.1         0.0001529 0.1        0.000153 0           0.0001539 0          0.000154 0.1         0.0001549 0.1        0.000155 0           0.0001559 0          0.000156 0           0.0001569 0          0.000157 0           0.0001579 0          0.000158 0.1         0.0001589 0.1        0.000159 0           0.0001599 0          0.00016 0.1          0.0001609 0.1        0.000161 0           0.0001619 0         )
Vcol_2 col_0_2 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0              6.9e-06 0            7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0            1.49e-05 0           1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0            2.29e-05 0           2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0              3.09e-05 0           3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.75         3.49e-05 0.75        3.5e-05 0            3.59e-05 0           3.6e-05 0.75         3.69e-05 0.75        3.7e-05 0            3.79e-05 0           3.8e-05 0            3.89e-05 0           3.9e-05 0            3.99e-05 0           4e-05 0.75           4.09e-05 0.75        4.1e-05 0            4.19e-05 0           4.2e-05 0.75         4.29e-05 0.75        4.3e-05 0            4.39e-05 0           4.4e-05 0.75         4.49e-05 0.75        4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 0.75         4.89e-05 0.75        4.9e-05 0            4.99e-05 0           5e-05 0.75           5.09e-05 0.75        5.1e-05 0            5.19e-05 0           5.2e-05 0.75         5.29e-05 0.75        5.3e-05 0            5.39e-05 0           5.4e-05 0            5.49e-05 0           5.5e-05 0            5.59e-05 0           5.6e-05 0.75         5.69e-05 0.75        5.7e-05 0            5.79e-05 0           5.8e-05 0.75         5.89e-05 0.75        5.9e-05 0            5.99e-05 0           6e-05 0.75           6.09e-05 0.75        6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 0.75         6.49e-05 0.75        6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0              7.09e-05 0           7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0            7.89e-05 0           7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0            8.69e-05 0           8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0            9.49e-05 0           9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.75         9.89e-05 0.75        9.9e-05 0            9.99e-05 0           0.0001 0.75          0.0001009 0.75       0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 0.75        0.0001049 0.75       0.000105 0           0.0001059 0          0.000106 0.75        0.0001069 0.75       0.000107 0           0.0001079 0          0.000108 0.75        0.0001089 0.75       0.000109 0           0.0001099 0          0.00011 0            0.0001109 0          0.000111 0           0.0001119 0          0.000112 0.75        0.0001129 0.75       0.000113 0           0.0001139 0          0.000114 0.75        0.0001149 0.75       0.000115 0           0.0001159 0          0.000116 0.75        0.0001169 0.75       0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 0.75         0.0001209 0.75       0.000121 0           0.0001219 0          0.000122 0.75        0.0001229 0.75       0.000123 0           0.0001239 0          0.000124 0.75        0.0001249 0.75       0.000125 0           0.0001259 0          0.000126 0           0.0001269 0          0.000127 0           0.0001279 0          0.000128 0.75        0.0001289 0.75       0.000129 0           0.0001299 0          0.00013 0.1          0.0001309 0.1        0.000131 0           0.0001319 0          0.000132 0.1         0.0001329 0.1        0.000133 0           0.0001339 0          0.000134 0           0.0001349 0          0.000135 0           0.0001359 0          0.000136 0.1         0.0001369 0.1        0.000137 0           0.0001379 0          0.000138 0.1         0.0001389 0.1        0.000139 0           0.0001399 0          0.00014 0.1          0.0001409 0.1        0.000141 0           0.0001419 0          0.000142 0           0.0001429 0          0.000143 0           0.0001439 0          0.000144 0.1         0.0001449 0.1        0.000145 0           0.0001459 0          0.000146 0.1         0.0001469 0.1        0.000147 0           0.0001479 0          0.000148 0.1         0.0001489 0.1        0.000149 0           0.0001499 0          0.00015 0            0.0001509 0          0.000151 0           0.0001519 0          0.000152 0.1         0.0001529 0.1        0.000153 0           0.0001539 0          0.000154 0.1         0.0001549 0.1        0.000155 0           0.0001559 0          0.000156 0.1         0.0001569 0.1        0.000157 0           0.0001579 0          0.000158 0           0.0001589 0          0.000159 0           0.0001599 0          0.00016 0.1          0.0001609 0.1        0.000161 0           0.0001619 0         )
Vcol_3 col_0_3 0 PWLZ(0 0                  9e-07 0              1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0              8.9e-06 0            9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0            1.69e-05 0           1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0            2.49e-05 0           2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0            3.29e-05 0           3.3e-05 0            3.39e-05 0           3.4e-05 0.75         3.49e-05 0.75        3.5e-05 0            3.59e-05 0           3.6e-05 0.75         3.69e-05 0.75        3.7e-05 0            3.79e-05 0           3.8e-05 0.75         3.89e-05 0.75        3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 0.75         4.29e-05 0.75        4.3e-05 0            4.39e-05 0           4.4e-05 0.75         4.49e-05 0.75        4.5e-05 0            4.59e-05 0           4.6e-05 0.75         4.69e-05 0.75        4.7e-05 0            4.79e-05 0           4.8e-05 0            4.89e-05 0           4.9e-05 0            4.99e-05 0           5e-05 0.75           5.09e-05 0.75        5.1e-05 0            5.19e-05 0           5.2e-05 0.75         5.29e-05 0.75        5.3e-05 0            5.39e-05 0           5.4e-05 0.75         5.49e-05 0.75        5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 0.75         5.89e-05 0.75        5.9e-05 0            5.99e-05 0           6e-05 0.75           6.09e-05 0.75        6.1e-05 0            6.19e-05 0           6.2e-05 0.75         6.29e-05 0.75        6.3e-05 0            6.39e-05 0           6.4e-05 0            6.49e-05 0           6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0            7.29e-05 0           7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0              8.09e-05 0           8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0            8.89e-05 0           8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0            9.69e-05 0           9.7e-05 0            9.79e-05 0           9.8e-05 0.75         9.89e-05 0.75        9.9e-05 0            9.99e-05 0           0.0001 0.75          0.0001009 0.75       0.000101 0           0.0001019 0          0.000102 0.75        0.0001029 0.75       0.000103 0           0.0001039 0          0.000104 0           0.0001049 0          0.000105 0           0.0001059 0          0.000106 0.75        0.0001069 0.75       0.000107 0           0.0001079 0          0.000108 0.75        0.0001089 0.75       0.000109 0           0.0001099 0          0.00011 0.75         0.0001109 0.75       0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 0.75        0.0001149 0.75       0.000115 0           0.0001159 0          0.000116 0.75        0.0001169 0.75       0.000117 0           0.0001179 0          0.000118 0.75        0.0001189 0.75       0.000119 0           0.0001199 0          0.00012 0            0.0001209 0          0.000121 0           0.0001219 0          0.000122 0.75        0.0001229 0.75       0.000123 0           0.0001239 0          0.000124 0.75        0.0001249 0.75       0.000125 0           0.0001259 0          0.000126 0.75        0.0001269 0.75       0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 0.1          0.0001309 0.1        0.000131 0           0.0001319 0          0.000132 0.1         0.0001329 0.1        0.000133 0           0.0001339 0          0.000134 0.1         0.0001349 0.1        0.000135 0           0.0001359 0          0.000136 0           0.0001369 0          0.000137 0           0.0001379 0          0.000138 0.1         0.0001389 0.1        0.000139 0           0.0001399 0          0.00014 0.1          0.0001409 0.1        0.000141 0           0.0001419 0          0.000142 0.1         0.0001429 0.1        0.000143 0           0.0001439 0          0.000144 0           0.0001449 0          0.000145 0           0.0001459 0          0.000146 0.1         0.0001469 0.1        0.000147 0           0.0001479 0          0.000148 0.1         0.0001489 0.1        0.000149 0           0.0001499 0          0.00015 0.1          0.0001509 0.1        0.000151 0           0.0001519 0          0.000152 0           0.0001529 0          0.000153 0           0.0001539 0          0.000154 0.1         0.0001549 0.1        0.000155 0           0.0001559 0          0.000156 0.1         0.0001569 0.1        0.000157 0           0.0001579 0          0.000158 0.1         0.0001589 0.1        0.000159 0           0.0001599 0          0.00016 0            0.0001609 0          0.000161 0           0.0001619 0         )


** Transient analysis **
.tran 1e-07 0.000162

.end