.title <test_2R_cb_8x8_2f>


** Includes **


** Load models **
.hdl ../models/rram_wp_akash.va

** Options **
.option post=2

** Parameters **


** Probes **


** Sub-circuits **
.subckt CELL r1 r2 c1 c2 mid gap1 gap2
Rr r1 r2 0.18
Cr r1 gnd 1.08e-13
Rc c1 c2 0.18
Cc c1 gnd 1.08e-13
X1 r1 mid gap1 RRAM_v0 
X2 c1 mid gap2 RRAM_v0 
.ends CELL


** Crossbar instantiation **
Xcell_0_0 row_0_0 row_0_1 col_0_0 col_1_0 mid_0_0 gap1_0_0 gap2_0_0 CELL
.ic v(gap1_0_0)=0.85 v(gap2_0_0)=0.85
Xcell_0_1 row_0_1 row_0_2 col_0_1 col_1_1 mid_0_1 gap1_0_1 gap2_0_1 CELL
.ic v(gap1_0_1)=0.85 v(gap2_0_1)=0.85
Xcell_0_2 row_0_2 row_0_3 col_0_2 col_1_2 mid_0_2 gap1_0_2 gap2_0_2 CELL
.ic v(gap1_0_2)=0.85 v(gap2_0_2)=0.85
Xcell_0_3 row_0_3 row_0_4 col_0_3 col_1_3 mid_0_3 gap1_0_3 gap2_0_3 CELL
.ic v(gap1_0_3)=0.85 v(gap2_0_3)=0.85
Xcell_0_4 row_0_4 row_0_5 col_0_4 col_1_4 mid_0_4 gap1_0_4 gap2_0_4 CELL
.ic v(gap1_0_4)=0.85 v(gap2_0_4)=0.85
Xcell_0_5 row_0_5 row_0_6 col_0_5 col_1_5 mid_0_5 gap1_0_5 gap2_0_5 CELL
.ic v(gap1_0_5)=0.85 v(gap2_0_5)=0.85
Xcell_0_6 row_0_6 row_0_7 col_0_6 col_1_6 mid_0_6 gap1_0_6 gap2_0_6 CELL
.ic v(gap1_0_6)=0.85 v(gap2_0_6)=0.85
Xcell_0_7 row_0_7 row_0_8 col_0_7 col_1_7 mid_0_7 gap1_0_7 gap2_0_7 CELL
.ic v(gap1_0_7)=0.85 v(gap2_0_7)=0.85
Xcell_1_0 row_1_0 row_1_1 col_1_0 col_2_0 mid_1_0 gap1_1_0 gap2_1_0 CELL
.ic v(gap1_1_0)=0.85 v(gap2_1_0)=0.85
Xcell_1_1 row_1_1 row_1_2 col_1_1 col_2_1 mid_1_1 gap1_1_1 gap2_1_1 CELL
.ic v(gap1_1_1)=0.85 v(gap2_1_1)=0.85
Xcell_1_2 row_1_2 row_1_3 col_1_2 col_2_2 mid_1_2 gap1_1_2 gap2_1_2 CELL
.ic v(gap1_1_2)=0.85 v(gap2_1_2)=0.85
Xcell_1_3 row_1_3 row_1_4 col_1_3 col_2_3 mid_1_3 gap1_1_3 gap2_1_3 CELL
.ic v(gap1_1_3)=0.85 v(gap2_1_3)=0.85
Xcell_1_4 row_1_4 row_1_5 col_1_4 col_2_4 mid_1_4 gap1_1_4 gap2_1_4 CELL
.ic v(gap1_1_4)=0.85 v(gap2_1_4)=0.85
Xcell_1_5 row_1_5 row_1_6 col_1_5 col_2_5 mid_1_5 gap1_1_5 gap2_1_5 CELL
.ic v(gap1_1_5)=0.85 v(gap2_1_5)=0.85
Xcell_1_6 row_1_6 row_1_7 col_1_6 col_2_6 mid_1_6 gap1_1_6 gap2_1_6 CELL
.ic v(gap1_1_6)=0.85 v(gap2_1_6)=0.85
Xcell_1_7 row_1_7 row_1_8 col_1_7 col_2_7 mid_1_7 gap1_1_7 gap2_1_7 CELL
.ic v(gap1_1_7)=0.85 v(gap2_1_7)=0.85
Xcell_2_0 row_2_0 row_2_1 col_2_0 col_3_0 mid_2_0 gap1_2_0 gap2_2_0 CELL
.ic v(gap1_2_0)=0.85 v(gap2_2_0)=0.85
Xcell_2_1 row_2_1 row_2_2 col_2_1 col_3_1 mid_2_1 gap1_2_1 gap2_2_1 CELL
.ic v(gap1_2_1)=0.85 v(gap2_2_1)=0.85
Xcell_2_2 row_2_2 row_2_3 col_2_2 col_3_2 mid_2_2 gap1_2_2 gap2_2_2 CELL
.ic v(gap1_2_2)=0.85 v(gap2_2_2)=0.85
Xcell_2_3 row_2_3 row_2_4 col_2_3 col_3_3 mid_2_3 gap1_2_3 gap2_2_3 CELL
.ic v(gap1_2_3)=0.85 v(gap2_2_3)=0.85
Xcell_2_4 row_2_4 row_2_5 col_2_4 col_3_4 mid_2_4 gap1_2_4 gap2_2_4 CELL
.ic v(gap1_2_4)=0.85 v(gap2_2_4)=0.85
Xcell_2_5 row_2_5 row_2_6 col_2_5 col_3_5 mid_2_5 gap1_2_5 gap2_2_5 CELL
.ic v(gap1_2_5)=0.85 v(gap2_2_5)=0.85
Xcell_2_6 row_2_6 row_2_7 col_2_6 col_3_6 mid_2_6 gap1_2_6 gap2_2_6 CELL
.ic v(gap1_2_6)=0.85 v(gap2_2_6)=0.85
Xcell_2_7 row_2_7 row_2_8 col_2_7 col_3_7 mid_2_7 gap1_2_7 gap2_2_7 CELL
.ic v(gap1_2_7)=0.85 v(gap2_2_7)=0.85
Xcell_3_0 row_3_0 row_3_1 col_3_0 col_4_0 mid_3_0 gap1_3_0 gap2_3_0 CELL
.ic v(gap1_3_0)=0.85 v(gap2_3_0)=0.85
Xcell_3_1 row_3_1 row_3_2 col_3_1 col_4_1 mid_3_1 gap1_3_1 gap2_3_1 CELL
.ic v(gap1_3_1)=0.85 v(gap2_3_1)=0.85
Xcell_3_2 row_3_2 row_3_3 col_3_2 col_4_2 mid_3_2 gap1_3_2 gap2_3_2 CELL
.ic v(gap1_3_2)=0.85 v(gap2_3_2)=0.85
Xcell_3_3 row_3_3 row_3_4 col_3_3 col_4_3 mid_3_3 gap1_3_3 gap2_3_3 CELL
.ic v(gap1_3_3)=0.85 v(gap2_3_3)=0.85
Xcell_3_4 row_3_4 row_3_5 col_3_4 col_4_4 mid_3_4 gap1_3_4 gap2_3_4 CELL
.ic v(gap1_3_4)=0.85 v(gap2_3_4)=0.85
Xcell_3_5 row_3_5 row_3_6 col_3_5 col_4_5 mid_3_5 gap1_3_5 gap2_3_5 CELL
.ic v(gap1_3_5)=0.85 v(gap2_3_5)=0.85
Xcell_3_6 row_3_6 row_3_7 col_3_6 col_4_6 mid_3_6 gap1_3_6 gap2_3_6 CELL
.ic v(gap1_3_6)=0.85 v(gap2_3_6)=0.85
Xcell_3_7 row_3_7 row_3_8 col_3_7 col_4_7 mid_3_7 gap1_3_7 gap2_3_7 CELL
.ic v(gap1_3_7)=0.85 v(gap2_3_7)=0.85
Xcell_4_0 row_4_0 row_4_1 col_4_0 col_5_0 mid_4_0 gap1_4_0 gap2_4_0 CELL
.ic v(gap1_4_0)=0.85 v(gap2_4_0)=0.85
Xcell_4_1 row_4_1 row_4_2 col_4_1 col_5_1 mid_4_1 gap1_4_1 gap2_4_1 CELL
.ic v(gap1_4_1)=0.85 v(gap2_4_1)=0.85
Xcell_4_2 row_4_2 row_4_3 col_4_2 col_5_2 mid_4_2 gap1_4_2 gap2_4_2 CELL
.ic v(gap1_4_2)=0.85 v(gap2_4_2)=0.85
Xcell_4_3 row_4_3 row_4_4 col_4_3 col_5_3 mid_4_3 gap1_4_3 gap2_4_3 CELL
.ic v(gap1_4_3)=0.85 v(gap2_4_3)=0.85
Xcell_4_4 row_4_4 row_4_5 col_4_4 col_5_4 mid_4_4 gap1_4_4 gap2_4_4 CELL
.ic v(gap1_4_4)=0.85 v(gap2_4_4)=0.85
Xcell_4_5 row_4_5 row_4_6 col_4_5 col_5_5 mid_4_5 gap1_4_5 gap2_4_5 CELL
.ic v(gap1_4_5)=0.85 v(gap2_4_5)=0.85
Xcell_4_6 row_4_6 row_4_7 col_4_6 col_5_6 mid_4_6 gap1_4_6 gap2_4_6 CELL
.ic v(gap1_4_6)=0.85 v(gap2_4_6)=0.85
Xcell_4_7 row_4_7 row_4_8 col_4_7 col_5_7 mid_4_7 gap1_4_7 gap2_4_7 CELL
.ic v(gap1_4_7)=0.85 v(gap2_4_7)=0.85
Xcell_5_0 row_5_0 row_5_1 col_5_0 col_6_0 mid_5_0 gap1_5_0 gap2_5_0 CELL
.ic v(gap1_5_0)=0.85 v(gap2_5_0)=0.85
Xcell_5_1 row_5_1 row_5_2 col_5_1 col_6_1 mid_5_1 gap1_5_1 gap2_5_1 CELL
.ic v(gap1_5_1)=0.85 v(gap2_5_1)=0.85
Xcell_5_2 row_5_2 row_5_3 col_5_2 col_6_2 mid_5_2 gap1_5_2 gap2_5_2 CELL
.ic v(gap1_5_2)=0.85 v(gap2_5_2)=0.85
Xcell_5_3 row_5_3 row_5_4 col_5_3 col_6_3 mid_5_3 gap1_5_3 gap2_5_3 CELL
.ic v(gap1_5_3)=0.85 v(gap2_5_3)=0.85
Xcell_5_4 row_5_4 row_5_5 col_5_4 col_6_4 mid_5_4 gap1_5_4 gap2_5_4 CELL
.ic v(gap1_5_4)=0.85 v(gap2_5_4)=0.85
Xcell_5_5 row_5_5 row_5_6 col_5_5 col_6_5 mid_5_5 gap1_5_5 gap2_5_5 CELL
.ic v(gap1_5_5)=0.85 v(gap2_5_5)=0.85
Xcell_5_6 row_5_6 row_5_7 col_5_6 col_6_6 mid_5_6 gap1_5_6 gap2_5_6 CELL
.ic v(gap1_5_6)=0.85 v(gap2_5_6)=0.85
Xcell_5_7 row_5_7 row_5_8 col_5_7 col_6_7 mid_5_7 gap1_5_7 gap2_5_7 CELL
.ic v(gap1_5_7)=0.85 v(gap2_5_7)=0.85
Xcell_6_0 row_6_0 row_6_1 col_6_0 col_7_0 mid_6_0 gap1_6_0 gap2_6_0 CELL
.ic v(gap1_6_0)=0.85 v(gap2_6_0)=0.85
Xcell_6_1 row_6_1 row_6_2 col_6_1 col_7_1 mid_6_1 gap1_6_1 gap2_6_1 CELL
.ic v(gap1_6_1)=0.85 v(gap2_6_1)=0.85
Xcell_6_2 row_6_2 row_6_3 col_6_2 col_7_2 mid_6_2 gap1_6_2 gap2_6_2 CELL
.ic v(gap1_6_2)=0.85 v(gap2_6_2)=0.85
Xcell_6_3 row_6_3 row_6_4 col_6_3 col_7_3 mid_6_3 gap1_6_3 gap2_6_3 CELL
.ic v(gap1_6_3)=0.85 v(gap2_6_3)=0.85
Xcell_6_4 row_6_4 row_6_5 col_6_4 col_7_4 mid_6_4 gap1_6_4 gap2_6_4 CELL
.ic v(gap1_6_4)=0.85 v(gap2_6_4)=0.85
Xcell_6_5 row_6_5 row_6_6 col_6_5 col_7_5 mid_6_5 gap1_6_5 gap2_6_5 CELL
.ic v(gap1_6_5)=0.85 v(gap2_6_5)=0.85
Xcell_6_6 row_6_6 row_6_7 col_6_6 col_7_6 mid_6_6 gap1_6_6 gap2_6_6 CELL
.ic v(gap1_6_6)=0.85 v(gap2_6_6)=0.85
Xcell_6_7 row_6_7 row_6_8 col_6_7 col_7_7 mid_6_7 gap1_6_7 gap2_6_7 CELL
.ic v(gap1_6_7)=0.85 v(gap2_6_7)=0.85
Xcell_7_0 row_7_0 row_7_1 col_7_0 col_8_0 mid_7_0 gap1_7_0 gap2_7_0 CELL
.ic v(gap1_7_0)=0.85 v(gap2_7_0)=0.85
Xcell_7_1 row_7_1 row_7_2 col_7_1 col_8_1 mid_7_1 gap1_7_1 gap2_7_1 CELL
.ic v(gap1_7_1)=0.85 v(gap2_7_1)=0.85
Xcell_7_2 row_7_2 row_7_3 col_7_2 col_8_2 mid_7_2 gap1_7_2 gap2_7_2 CELL
.ic v(gap1_7_2)=0.85 v(gap2_7_2)=0.85
Xcell_7_3 row_7_3 row_7_4 col_7_3 col_8_3 mid_7_3 gap1_7_3 gap2_7_3 CELL
.ic v(gap1_7_3)=0.85 v(gap2_7_3)=0.85
Xcell_7_4 row_7_4 row_7_5 col_7_4 col_8_4 mid_7_4 gap1_7_4 gap2_7_4 CELL
.ic v(gap1_7_4)=0.85 v(gap2_7_4)=0.85
Xcell_7_5 row_7_5 row_7_6 col_7_5 col_8_5 mid_7_5 gap1_7_5 gap2_7_5 CELL
.ic v(gap1_7_5)=0.85 v(gap2_7_5)=0.85
Xcell_7_6 row_7_6 row_7_7 col_7_6 col_8_6 mid_7_6 gap1_7_6 gap2_7_6 CELL
.ic v(gap1_7_6)=0.85 v(gap2_7_6)=0.85
Xcell_7_7 row_7_7 row_7_8 col_7_7 col_8_7 mid_7_7 gap1_7_7 gap2_7_7 CELL
.ic v(gap1_7_7)=0.85 v(gap2_7_7)=0.85


** PWL voltage waveforms **
Vrow_0 row_0_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 3              4.9e-06 3            5e-06 0              5.9e-06 0            6e-06 0              6.9e-06 0            7e-06 0              7.9e-06 0            8e-06 3              8.9e-06 3            9e-06 0              9.9e-06 0            1e-05 0              1.09e-05 0           1.1e-05 0            1.19e-05 0           1.2e-05 3            1.29e-05 3           1.3e-05 0            1.39e-05 0           1.4e-05 0            1.49e-05 0           1.5e-05 0            1.59e-05 0           1.6e-05 3            1.69e-05 3           1.7e-05 0            1.79e-05 0           1.8e-05 0            1.89e-05 0           1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 0           0.0001349 0          0.000135 0           0.0001359 0          0.000136 3           0.0001369 3          0.000137 0           0.0001379 0          0.000138 0           0.0001389 0          0.000139 0           0.0001399 0          0.00014 3            0.0001409 3          0.000141 0           0.0001419 0          0.000142 0           0.0001429 0          0.000143 0           0.0001439 0          0.000144 3           0.0001449 3          0.000145 0           0.0001459 0          0.000146 0           0.0001469 0          0.000147 0           0.0001479 0          0.000148 3           0.0001489 3          0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_1 row_1_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 0              2.09e-05 0           2.1e-05 0            2.19e-05 0           2.2e-05 3            2.29e-05 3           2.3e-05 0            2.39e-05 0           2.4e-05 0            2.49e-05 0           2.5e-05 0            2.59e-05 0           2.6e-05 3            2.69e-05 3           2.7e-05 0            2.79e-05 0           2.8e-05 0            2.89e-05 0           2.9e-05 0            2.99e-05 0           3e-05 3              3.09e-05 3           3.1e-05 0            3.19e-05 0           3.2e-05 0            3.29e-05 0           3.3e-05 0            3.39e-05 0           3.4e-05 3            3.49e-05 3           3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 3            0.0001509 3          0.000151 0           0.0001519 0          0.000152 0           0.0001529 0          0.000153 0           0.0001539 0          0.000154 3           0.0001549 3          0.000155 0           0.0001559 0          0.000156 0           0.0001569 0          0.000157 0           0.0001579 0          0.000158 3           0.0001589 3          0.000159 0           0.0001599 0          0.00016 0            0.0001609 0          0.000161 0           0.0001619 0          0.000162 3           0.0001629 3          0.000163 0           0.0001639 0          0.000164 0           0.0001649 0          0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_2 row_2_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 3            3.69e-05 3           3.7e-05 0            3.79e-05 0           3.8e-05 0            3.89e-05 0           3.9e-05 0            3.99e-05 0           4e-05 3              4.09e-05 3           4.1e-05 0            4.19e-05 0           4.2e-05 0            4.29e-05 0           4.3e-05 0            4.39e-05 0           4.4e-05 3            4.49e-05 3           4.5e-05 0            4.59e-05 0           4.6e-05 0            4.69e-05 0           4.7e-05 0            4.79e-05 0           4.8e-05 3            4.89e-05 3           4.9e-05 0            4.99e-05 0           5e-05 0              5.09e-05 0           5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 0           0.0001669 0          0.000167 0           0.0001679 0          0.000168 3           0.0001689 3          0.000169 0           0.0001699 0          0.00017 0            0.0001709 0          0.000171 0           0.0001719 0          0.000172 3           0.0001729 3          0.000173 0           0.0001739 0          0.000174 0           0.0001749 0          0.000175 0           0.0001759 0          0.000176 3           0.0001769 3          0.000177 0           0.0001779 0          0.000178 0           0.0001789 0          0.000179 0           0.0001799 0          0.00018 3            0.0001809 3          0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_3 row_3_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 0            5.29e-05 0           5.3e-05 0            5.39e-05 0           5.4e-05 3            5.49e-05 3           5.5e-05 0            5.59e-05 0           5.6e-05 0            5.69e-05 0           5.7e-05 0            5.79e-05 0           5.8e-05 3            5.89e-05 3           5.9e-05 0            5.99e-05 0           6e-05 0              6.09e-05 0           6.1e-05 0            6.19e-05 0           6.2e-05 3            6.29e-05 3           6.3e-05 0            6.39e-05 0           6.4e-05 0            6.49e-05 0           6.5e-05 0            6.59e-05 0           6.6e-05 3            6.69e-05 3           6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 3           0.0001829 3          0.000183 0           0.0001839 0          0.000184 0           0.0001849 0          0.000185 0           0.0001859 0          0.000186 3           0.0001869 3          0.000187 0           0.0001879 0          0.000188 0           0.0001889 0          0.000189 0           0.0001899 0          0.00019 3            0.0001909 3          0.000191 0           0.0001919 0          0.000192 0           0.0001929 0          0.000193 0           0.0001939 0          0.000194 3           0.0001949 3          0.000195 0           0.0001959 0          0.000196 0           0.0001969 0          0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_4 row_4_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 3            6.89e-05 3           6.9e-05 0            6.99e-05 0           7e-05 0              7.09e-05 0           7.1e-05 0            7.19e-05 0           7.2e-05 3            7.29e-05 3           7.3e-05 0            7.39e-05 0           7.4e-05 0            7.49e-05 0           7.5e-05 0            7.59e-05 0           7.6e-05 3            7.69e-05 3           7.7e-05 0            7.79e-05 0           7.8e-05 0            7.89e-05 0           7.9e-05 0            7.99e-05 0           8e-05 3              8.09e-05 3           8.1e-05 0            8.19e-05 0           8.2e-05 0            8.29e-05 0           8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 0           0.0001989 0          0.000199 0           0.0001999 0          0.0002 3             0.0002009 3          0.000201 0           0.0002019 0          0.000202 0           0.0002029 0          0.000203 0           0.0002039 0          0.000204 3           0.0002049 3          0.000205 0           0.0002059 0          0.000206 0           0.0002069 0          0.000207 0           0.0002079 0          0.000208 3           0.0002089 3          0.000209 0           0.0002099 0          0.00021 0            0.0002109 0          0.000211 0           0.0002119 0          0.000212 3           0.0002129 3          0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_5 row_5_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 0            8.49e-05 0           8.5e-05 0            8.59e-05 0           8.6e-05 3            8.69e-05 3           8.7e-05 0            8.79e-05 0           8.8e-05 0            8.89e-05 0           8.9e-05 0            8.99e-05 0           9e-05 3              9.09e-05 3           9.1e-05 0            9.19e-05 0           9.2e-05 0            9.29e-05 0           9.3e-05 0            9.39e-05 0           9.4e-05 3            9.49e-05 3           9.5e-05 0            9.59e-05 0           9.6e-05 0            9.69e-05 0           9.7e-05 0            9.79e-05 0           9.8e-05 3            9.89e-05 3           9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 3           0.0002149 3          0.000215 0           0.0002159 0          0.000216 0           0.0002169 0          0.000217 0           0.0002179 0          0.000218 3           0.0002189 3          0.000219 0           0.0002199 0          0.00022 0            0.0002209 0          0.000221 0           0.0002219 0          0.000222 3           0.0002229 3          0.000223 0           0.0002239 0          0.000224 0           0.0002249 0          0.000225 0           0.0002259 0          0.000226 3           0.0002269 3          0.000227 0           0.0002279 0          0.000228 0           0.0002289 0          0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_6 row_6_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 3             0.0001009 3          0.000101 0           0.0001019 0          0.000102 0           0.0001029 0          0.000103 0           0.0001039 0          0.000104 3           0.0001049 3          0.000105 0           0.0001059 0          0.000106 0           0.0001069 0          0.000107 0           0.0001079 0          0.000108 3           0.0001089 3          0.000109 0           0.0001099 0          0.00011 0            0.0001109 0          0.000111 0           0.0001119 0          0.000112 3           0.0001129 3          0.000113 0           0.0001139 0          0.000114 0           0.0001149 0          0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 0            0.0002309 0          0.000231 0           0.0002319 0          0.000232 3           0.0002329 3          0.000233 0           0.0002339 0          0.000234 0           0.0002349 0          0.000235 0           0.0002359 0          0.000236 3           0.0002369 3          0.000237 0           0.0002379 0          0.000238 0           0.0002389 0          0.000239 0           0.0002399 0          0.00024 3            0.0002409 3          0.000241 0           0.0002419 0          0.000242 0           0.0002429 0          0.000243 0           0.0002439 0          0.000244 3           0.0002449 3          0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vrow_7 row_7_0 0 PWLZ(0 0                  9e-07 0              1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 0           0.0001169 0          0.000117 0           0.0001179 0          0.000118 3           0.0001189 3          0.000119 0           0.0001199 0          0.00012 0            0.0001209 0          0.000121 0           0.0001219 0          0.000122 3           0.0001229 3          0.000123 0           0.0001239 0          0.000124 0           0.0001249 0          0.000125 0           0.0001259 0          0.000126 3           0.0001269 3          0.000127 0           0.0001279 0          0.000128 0           0.0001289 0          0.000129 0           0.0001299 0          0.00013 3            0.0001309 3          0.000131 0           0.0001319 0          0.000132 0.2         0.0001329 0.2        0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 3           0.0002469 3          0.000247 0           0.0002479 0          0.000248 0           0.0002489 0          0.000249 0           0.0002499 0          0.00025 3            0.0002509 3          0.000251 0           0.0002519 0          0.000252 0           0.0002529 0          0.000253 0           0.0002539 0          0.000254 3           0.0002549 3          0.000255 0           0.0002559 0          0.000256 0           0.0002569 0          0.000257 0           0.0002579 0          0.000258 3           0.0002589 3          0.000259 0           0.0002599 0          0.00026 0            0.0002609 0          0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0         )
Vcol_0 col_0_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 0              4.9e-06 0            5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 3              2.09e-05 3           2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 0            3.69e-05 0           3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 3            5.29e-05 3           5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 0            6.89e-05 0           6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 3            8.49e-05 3           8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 0             0.0001009 0          0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 3           0.0001169 3          0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 3           0.0001349 3          0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 0            0.0001509 0          0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 3           0.0001669 3          0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 0           0.0001829 0          0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 3           0.0001989 3          0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 0           0.0002149 0          0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 3            0.0002309 3          0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 0           0.0002469 0          0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_1 col_0_1 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 3              6.9e-06 3            7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 0            2.29e-05 0           2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 3            3.89e-05 3           3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 0            5.49e-05 0           5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 3              7.09e-05 3           7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 0            8.69e-05 0           8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 3           0.0001029 3          0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 0           0.0001189 0          0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 0           0.0001369 0          0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 3           0.0001529 3          0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 0           0.0001689 0          0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 3           0.0001849 3          0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 0             0.0002009 0          0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 3           0.0002169 3          0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 0           0.0002329 0          0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 3           0.0002489 3          0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_2 col_0_2 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 0              8.9e-06 0            9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 3            2.49e-05 3           2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 0              4.09e-05 0           4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 3            5.69e-05 3           5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 0            7.29e-05 0           7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 3            8.89e-05 3           8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 0           0.0001049 0          0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 3            0.0001209 3          0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 3           0.0001389 3          0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 0           0.0001549 0          0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 3            0.0001709 3          0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 0           0.0001869 0          0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 3           0.0002029 3          0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 0           0.0002189 0          0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 3           0.0002349 3          0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 0            0.0002509 0          0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_3 col_0_3 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 3              1.09e-05 3           1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 0            2.69e-05 0           2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 3            4.29e-05 3           4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 0            5.89e-05 0           5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 3            7.49e-05 3           7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 0              9.09e-05 0           9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 3           0.0001069 3          0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 0           0.0001229 0          0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 0            0.0001409 0          0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 3           0.0001569 3          0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 0           0.0001729 0          0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 3           0.0001889 3          0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 0           0.0002049 0          0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 3            0.0002209 3          0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 0           0.0002369 0          0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 3           0.0002529 3          0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_4 col_0_4 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 0            1.29e-05 0           1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 3            2.89e-05 3           2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 0            4.49e-05 0           4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 3              6.09e-05 3           6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 0            7.69e-05 0           7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 3            9.29e-05 3           9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 0           0.0001089 0          0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 3           0.0001249 3          0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 3           0.0001429 3          0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 0           0.0001589 0          0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 3           0.0001749 3          0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 0            0.0001909 0          0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 3           0.0002069 3          0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 0           0.0002229 0          0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 3           0.0002389 3          0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 0           0.0002549 0          0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_5 col_0_5 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 3            1.49e-05 3           1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 0              3.09e-05 0           3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 3            4.69e-05 3           4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 0            6.29e-05 0           6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 3            7.89e-05 3           7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 0            9.49e-05 0           9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 3            0.0001109 3          0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 0           0.0001269 0          0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 0           0.0001449 0          0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 3            0.0001609 3          0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 0           0.0001769 0          0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 3           0.0001929 3          0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 0           0.0002089 0          0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 3           0.0002249 3          0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 0            0.0002409 0          0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 3           0.0002569 3          0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_6 col_0_6 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 0            1.69e-05 0           1.7e-05 0            1.79e-05 0           1.8e-05 1.5          1.89e-05 1.5         1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 3            3.29e-05 3           3.3e-05 0            3.39e-05 0           3.4e-05 1.5          3.49e-05 1.5         3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 0            4.89e-05 0           4.9e-05 0            4.99e-05 0           5e-05 1.5            5.09e-05 1.5         5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 3            6.49e-05 3           6.5e-05 0            6.59e-05 0           6.6e-05 1.5          6.69e-05 1.5         6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 0              8.09e-05 0           8.1e-05 0            8.19e-05 0           8.2e-05 1.5          8.29e-05 1.5         8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 3            9.69e-05 3           9.7e-05 0            9.79e-05 0           9.8e-05 1.5          9.89e-05 1.5         9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 0           0.0001129 0          0.000113 0           0.0001139 0          0.000114 1.5         0.0001149 1.5        0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 3           0.0001289 3          0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 3           0.0001469 3          0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 0           0.0001629 0          0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 3           0.0001789 3          0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 0           0.0001949 0          0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 3            0.0002109 3          0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 0           0.0002269 0          0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 3           0.0002429 3          0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 0           0.0002589 0          0.000259 0           0.0002599 0          0.00026 1.5          0.0002609 1.5        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )
Vcol_7 col_0_7 0 PWLZ(0 0                  9e-07 0              1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 1.5            4.9e-06 1.5          5e-06 0              5.9e-06 0            6e-06 1.5            6.9e-06 1.5          7e-06 0              7.9e-06 0            8e-06 1.5            8.9e-06 1.5          9e-06 0              9.9e-06 0            1e-05 1.5            1.09e-05 1.5         1.1e-05 0            1.19e-05 0           1.2e-05 1.5          1.29e-05 1.5         1.3e-05 0            1.39e-05 0           1.4e-05 1.5          1.49e-05 1.5         1.5e-05 0            1.59e-05 0           1.6e-05 1.5          1.69e-05 1.5         1.7e-05 0            1.79e-05 0           1.8e-05 3            1.89e-05 3           1.9e-05 0            1.99e-05 0           2e-05 1.5            2.09e-05 1.5         2.1e-05 0            2.19e-05 0           2.2e-05 1.5          2.29e-05 1.5         2.3e-05 0            2.39e-05 0           2.4e-05 1.5          2.49e-05 1.5         2.5e-05 0            2.59e-05 0           2.6e-05 1.5          2.69e-05 1.5         2.7e-05 0            2.79e-05 0           2.8e-05 1.5          2.89e-05 1.5         2.9e-05 0            2.99e-05 0           3e-05 1.5            3.09e-05 1.5         3.1e-05 0            3.19e-05 0           3.2e-05 1.5          3.29e-05 1.5         3.3e-05 0            3.39e-05 0           3.4e-05 0            3.49e-05 0           3.5e-05 0            3.59e-05 0           3.6e-05 1.5          3.69e-05 1.5         3.7e-05 0            3.79e-05 0           3.8e-05 1.5          3.89e-05 1.5         3.9e-05 0            3.99e-05 0           4e-05 1.5            4.09e-05 1.5         4.1e-05 0            4.19e-05 0           4.2e-05 1.5          4.29e-05 1.5         4.3e-05 0            4.39e-05 0           4.4e-05 1.5          4.49e-05 1.5         4.5e-05 0            4.59e-05 0           4.6e-05 1.5          4.69e-05 1.5         4.7e-05 0            4.79e-05 0           4.8e-05 1.5          4.89e-05 1.5         4.9e-05 0            4.99e-05 0           5e-05 3              5.09e-05 3           5.1e-05 0            5.19e-05 0           5.2e-05 1.5          5.29e-05 1.5         5.3e-05 0            5.39e-05 0           5.4e-05 1.5          5.49e-05 1.5         5.5e-05 0            5.59e-05 0           5.6e-05 1.5          5.69e-05 1.5         5.7e-05 0            5.79e-05 0           5.8e-05 1.5          5.89e-05 1.5         5.9e-05 0            5.99e-05 0           6e-05 1.5            6.09e-05 1.5         6.1e-05 0            6.19e-05 0           6.2e-05 1.5          6.29e-05 1.5         6.3e-05 0            6.39e-05 0           6.4e-05 1.5          6.49e-05 1.5         6.5e-05 0            6.59e-05 0           6.6e-05 0            6.69e-05 0           6.7e-05 0            6.79e-05 0           6.8e-05 1.5          6.89e-05 1.5         6.9e-05 0            6.99e-05 0           7e-05 1.5            7.09e-05 1.5         7.1e-05 0            7.19e-05 0           7.2e-05 1.5          7.29e-05 1.5         7.3e-05 0            7.39e-05 0           7.4e-05 1.5          7.49e-05 1.5         7.5e-05 0            7.59e-05 0           7.6e-05 1.5          7.69e-05 1.5         7.7e-05 0            7.79e-05 0           7.8e-05 1.5          7.89e-05 1.5         7.9e-05 0            7.99e-05 0           8e-05 1.5            8.09e-05 1.5         8.1e-05 0            8.19e-05 0           8.2e-05 3            8.29e-05 3           8.3e-05 0            8.39e-05 0           8.4e-05 1.5          8.49e-05 1.5         8.5e-05 0            8.59e-05 0           8.6e-05 1.5          8.69e-05 1.5         8.7e-05 0            8.79e-05 0           8.8e-05 1.5          8.89e-05 1.5         8.9e-05 0            8.99e-05 0           9e-05 1.5            9.09e-05 1.5         9.1e-05 0            9.19e-05 0           9.2e-05 1.5          9.29e-05 1.5         9.3e-05 0            9.39e-05 0           9.4e-05 1.5          9.49e-05 1.5         9.5e-05 0            9.59e-05 0           9.6e-05 1.5          9.69e-05 1.5         9.7e-05 0            9.79e-05 0           9.8e-05 0            9.89e-05 0           9.9e-05 0            9.99e-05 0           0.0001 1.5           0.0001009 1.5        0.000101 0           0.0001019 0          0.000102 1.5         0.0001029 1.5        0.000103 0           0.0001039 0          0.000104 1.5         0.0001049 1.5        0.000105 0           0.0001059 0          0.000106 1.5         0.0001069 1.5        0.000107 0           0.0001079 0          0.000108 1.5         0.0001089 1.5        0.000109 0           0.0001099 0          0.00011 1.5          0.0001109 1.5        0.000111 0           0.0001119 0          0.000112 1.5         0.0001129 1.5        0.000113 0           0.0001139 0          0.000114 3           0.0001149 3          0.000115 0           0.0001159 0          0.000116 1.5         0.0001169 1.5        0.000117 0           0.0001179 0          0.000118 1.5         0.0001189 1.5        0.000119 0           0.0001199 0          0.00012 1.5          0.0001209 1.5        0.000121 0           0.0001219 0          0.000122 1.5         0.0001229 1.5        0.000123 0           0.0001239 0          0.000124 1.5         0.0001249 1.5        0.000125 0           0.0001259 0          0.000126 1.5         0.0001269 1.5        0.000127 0           0.0001279 0          0.000128 1.5         0.0001289 1.5        0.000129 0           0.0001299 0          0.00013 0            0.0001309 0          0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 0           0.0001489 0          0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 3           0.0001649 3          0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 0            0.0001809 0          0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 3           0.0001969 3          0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 0           0.0002129 0          0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 3           0.0002289 3          0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 0           0.0002449 0          0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 1.5         0.0002589 1.5        0.000259 0           0.0002599 0          0.00026 3            0.0002609 3          0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0         )


** Transient analysis **
.tran 1e-07 0.000264

.end