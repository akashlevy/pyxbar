.title <test_1R_cb_8x8_2f>


** Includes **


** Load models **
.hdl ../models/rram_wp.va

** Options **
.option post=2

** Parameters **


** Probes **


** Sub-circuits **
.subckt CELL r1 r2 c1 c2 gap
Rr r1 r2 0.18
Cr r2 gnd 1.08e-13
Rc c1 c2 0.18
Cc c2 gnd 1.08e-13
X1 r1 c1 gap RRAM_v0 
.ends CELL


** Crossbar instantiation **
Xcell_0_0 row_0_0 row_0_1 col_0_0 col_1_0 gap_0_0 CELL
Xcell_0_1 row_0_1 row_0_2 col_0_1 col_1_1 gap_0_1 CELL
Xcell_0_2 row_0_2 row_0_3 col_0_2 col_1_2 gap_0_2 CELL
Xcell_0_3 row_0_3 row_0_4 col_0_3 col_1_3 gap_0_3 CELL
Xcell_0_4 row_0_4 row_0_5 col_0_4 col_1_4 gap_0_4 CELL
Xcell_0_5 row_0_5 row_0_6 col_0_5 col_1_5 gap_0_5 CELL
Xcell_0_6 row_0_6 row_0_7 col_0_6 col_1_6 gap_0_6 CELL
Xcell_0_7 row_0_7 row_0_8 col_0_7 col_1_7 gap_0_7 CELL
Xcell_1_0 row_1_0 row_1_1 col_1_0 col_2_0 gap_1_0 CELL
Xcell_1_1 row_1_1 row_1_2 col_1_1 col_2_1 gap_1_1 CELL
Xcell_1_2 row_1_2 row_1_3 col_1_2 col_2_2 gap_1_2 CELL
Xcell_1_3 row_1_3 row_1_4 col_1_3 col_2_3 gap_1_3 CELL
Xcell_1_4 row_1_4 row_1_5 col_1_4 col_2_4 gap_1_4 CELL
Xcell_1_5 row_1_5 row_1_6 col_1_5 col_2_5 gap_1_5 CELL
Xcell_1_6 row_1_6 row_1_7 col_1_6 col_2_6 gap_1_6 CELL
Xcell_1_7 row_1_7 row_1_8 col_1_7 col_2_7 gap_1_7 CELL
Xcell_2_0 row_2_0 row_2_1 col_2_0 col_3_0 gap_2_0 CELL
Xcell_2_1 row_2_1 row_2_2 col_2_1 col_3_1 gap_2_1 CELL
Xcell_2_2 row_2_2 row_2_3 col_2_2 col_3_2 gap_2_2 CELL
Xcell_2_3 row_2_3 row_2_4 col_2_3 col_3_3 gap_2_3 CELL
Xcell_2_4 row_2_4 row_2_5 col_2_4 col_3_4 gap_2_4 CELL
Xcell_2_5 row_2_5 row_2_6 col_2_5 col_3_5 gap_2_5 CELL
Xcell_2_6 row_2_6 row_2_7 col_2_6 col_3_6 gap_2_6 CELL
Xcell_2_7 row_2_7 row_2_8 col_2_7 col_3_7 gap_2_7 CELL
Xcell_3_0 row_3_0 row_3_1 col_3_0 col_4_0 gap_3_0 CELL
Xcell_3_1 row_3_1 row_3_2 col_3_1 col_4_1 gap_3_1 CELL
Xcell_3_2 row_3_2 row_3_3 col_3_2 col_4_2 gap_3_2 CELL
Xcell_3_3 row_3_3 row_3_4 col_3_3 col_4_3 gap_3_3 CELL
Xcell_3_4 row_3_4 row_3_5 col_3_4 col_4_4 gap_3_4 CELL
Xcell_3_5 row_3_5 row_3_6 col_3_5 col_4_5 gap_3_5 CELL
Xcell_3_6 row_3_6 row_3_7 col_3_6 col_4_6 gap_3_6 CELL
Xcell_3_7 row_3_7 row_3_8 col_3_7 col_4_7 gap_3_7 CELL
Xcell_4_0 row_4_0 row_4_1 col_4_0 col_5_0 gap_4_0 CELL
Xcell_4_1 row_4_1 row_4_2 col_4_1 col_5_1 gap_4_1 CELL
Xcell_4_2 row_4_2 row_4_3 col_4_2 col_5_2 gap_4_2 CELL
Xcell_4_3 row_4_3 row_4_4 col_4_3 col_5_3 gap_4_3 CELL
Xcell_4_4 row_4_4 row_4_5 col_4_4 col_5_4 gap_4_4 CELL
Xcell_4_5 row_4_5 row_4_6 col_4_5 col_5_5 gap_4_5 CELL
Xcell_4_6 row_4_6 row_4_7 col_4_6 col_5_6 gap_4_6 CELL
Xcell_4_7 row_4_7 row_4_8 col_4_7 col_5_7 gap_4_7 CELL
Xcell_5_0 row_5_0 row_5_1 col_5_0 col_6_0 gap_5_0 CELL
Xcell_5_1 row_5_1 row_5_2 col_5_1 col_6_1 gap_5_1 CELL
Xcell_5_2 row_5_2 row_5_3 col_5_2 col_6_2 gap_5_2 CELL
Xcell_5_3 row_5_3 row_5_4 col_5_3 col_6_3 gap_5_3 CELL
Xcell_5_4 row_5_4 row_5_5 col_5_4 col_6_4 gap_5_4 CELL
Xcell_5_5 row_5_5 row_5_6 col_5_5 col_6_5 gap_5_5 CELL
Xcell_5_6 row_5_6 row_5_7 col_5_6 col_6_6 gap_5_6 CELL
Xcell_5_7 row_5_7 row_5_8 col_5_7 col_6_7 gap_5_7 CELL
Xcell_6_0 row_6_0 row_6_1 col_6_0 col_7_0 gap_6_0 CELL
Xcell_6_1 row_6_1 row_6_2 col_6_1 col_7_1 gap_6_1 CELL
Xcell_6_2 row_6_2 row_6_3 col_6_2 col_7_2 gap_6_2 CELL
Xcell_6_3 row_6_3 row_6_4 col_6_3 col_7_3 gap_6_3 CELL
Xcell_6_4 row_6_4 row_6_5 col_6_4 col_7_4 gap_6_4 CELL
Xcell_6_5 row_6_5 row_6_6 col_6_5 col_7_5 gap_6_5 CELL
Xcell_6_6 row_6_6 row_6_7 col_6_6 col_7_6 gap_6_6 CELL
Xcell_6_7 row_6_7 row_6_8 col_6_7 col_7_7 gap_6_7 CELL
Xcell_7_0 row_7_0 row_7_1 col_7_0 col_8_0 gap_7_0 CELL
Xcell_7_1 row_7_1 row_7_2 col_7_1 col_8_1 gap_7_1 CELL
Xcell_7_2 row_7_2 row_7_3 col_7_2 col_8_2 gap_7_2 CELL
Xcell_7_3 row_7_3 row_7_4 col_7_3 col_8_3 gap_7_3 CELL
Xcell_7_4 row_7_4 row_7_5 col_7_4 col_8_4 gap_7_4 CELL
Xcell_7_5 row_7_5 row_7_6 col_7_5 col_8_5 gap_7_5 CELL
Xcell_7_6 row_7_6 row_7_7 col_7_6 col_8_6 gap_7_6 CELL
Xcell_7_7 row_7_7 row_7_8 col_7_7 col_8_7 gap_7_7 CELL


** PWL voltage waveforms **
Vrow_0 row_0_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.2            2.9e-06 0.2          3e-06 0              3.9e-06 0            4e-06 0.2            4.9e-06 0.2          5e-06 0              5.9e-06 0            6e-06 0.2            6.9e-06 0.2          7e-06 0              7.9e-06 0            8e-06 0.2            8.9e-06 0.2          9e-06 0              9.9e-06 0            1e-05 0.2            1.09e-05 0.2         1.1e-05 0            1.19e-05 0           1.2e-05 0.2          1.29e-05 0.2         1.3e-05 0            1.39e-05 0           1.4e-05 0.2          1.49e-05 0.2         1.5e-05 0            1.59e-05 0           1.6e-05 0.2          1.69e-05 0.2         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 1.5          0.0001309 1.5        0.000131 0           0.0001319 0          0.000132 0           0.0001329 0          0.000133 0           0.0001339 0          0.000134 1.5         0.0001349 1.5        0.000135 0           0.0001359 0          0.000136 0           0.0001369 0          0.000137 0           0.0001379 0          0.000138 1.5         0.0001389 1.5        0.000139 0           0.0001399 0          0.00014 0            0.0001409 0          0.000141 0           0.0001419 0          0.000142 1.5         0.0001429 1.5        0.000143 0           0.0001439 0          0.000144 0           0.0001449 0          0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.2         0.0002589 0.2        0.000259 0           0.0002599 0          0.00026 0.2          0.0002609 0.2        0.000261 0           0.0002619 0          0.000262 0.2         0.0002629 0.2        0.000263 0           0.0002639 0          0.000264 0.2         0.0002649 0.2        0.000265 0           0.0002659 0          0.000266 0.2         0.0002669 0.2        0.000267 0           0.0002679 0          0.000268 0.2         0.0002689 0.2        0.000269 0           0.0002699 0          0.00027 0.2          0.0002709 0.2        0.000271 0           0.0002719 0          0.000272 0.2         0.0002729 0.2        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0           0.0003869 0          0.000387 0           0.0003879 0          0.000388 1.5         0.0003889 1.5        0.000389 0           0.0003899 0          0.00039 0            0.0003909 0          0.000391 0           0.0003919 0          0.000392 1.5         0.0003929 1.5        0.000393 0           0.0003939 0          0.000394 0           0.0003949 0          0.000395 0           0.0003959 0          0.000396 1.5         0.0003969 1.5        0.000397 0           0.0003979 0          0.000398 0           0.0003989 0          0.000399 0           0.0003999 0          0.0004 1.5           0.0004009 1.5        0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.2         0.0005149 0.2        0.000515 0           0.0005159 0          0.000516 0.2         0.0005169 0.2        0.000517 0           0.0005179 0          0.000518 0.2         0.0005189 0.2        0.000519 0           0.0005199 0          0.00052 0.2          0.0005209 0.2        0.000521 0           0.0005219 0          0.000522 0.2         0.0005229 0.2        0.000523 0           0.0005239 0          0.000524 0.2         0.0005249 0.2        0.000525 0           0.0005259 0          0.000526 0.2         0.0005269 0.2        0.000527 0           0.0005279 0          0.000528 0.2         0.0005289 0.2        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_1 row_1_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.2          1.89e-05 0.2         1.9e-05 0            1.99e-05 0           2e-05 0.2            2.09e-05 0.2         2.1e-05 0            2.19e-05 0           2.2e-05 0.2          2.29e-05 0.2         2.3e-05 0            2.39e-05 0           2.4e-05 0.2          2.49e-05 0.2         2.5e-05 0            2.59e-05 0           2.6e-05 0.2          2.69e-05 0.2         2.7e-05 0            2.79e-05 0           2.8e-05 0.2          2.89e-05 0.2         2.9e-05 0            2.99e-05 0           3e-05 0.2            3.09e-05 0.2         3.1e-05 0            3.19e-05 0           3.2e-05 0.2          3.29e-05 0.2         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0           0.0001469 0          0.000147 0           0.0001479 0          0.000148 1.5         0.0001489 1.5        0.000149 0           0.0001499 0          0.00015 0            0.0001509 0          0.000151 0           0.0001519 0          0.000152 1.5         0.0001529 1.5        0.000153 0           0.0001539 0          0.000154 0           0.0001549 0          0.000155 0           0.0001559 0          0.000156 1.5         0.0001569 1.5        0.000157 0           0.0001579 0          0.000158 0           0.0001589 0          0.000159 0           0.0001599 0          0.00016 1.5          0.0001609 1.5        0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.2         0.0002749 0.2        0.000275 0           0.0002759 0          0.000276 0.2         0.0002769 0.2        0.000277 0           0.0002779 0          0.000278 0.2         0.0002789 0.2        0.000279 0           0.0002799 0          0.00028 0.2          0.0002809 0.2        0.000281 0           0.0002819 0          0.000282 0.2         0.0002829 0.2        0.000283 0           0.0002839 0          0.000284 0.2         0.0002849 0.2        0.000285 0           0.0002859 0          0.000286 0.2         0.0002869 0.2        0.000287 0           0.0002879 0          0.000288 0.2         0.0002889 0.2        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 1.5         0.0004029 1.5        0.000403 0           0.0004039 0          0.000404 0           0.0004049 0          0.000405 0           0.0004059 0          0.000406 1.5         0.0004069 1.5        0.000407 0           0.0004079 0          0.000408 0           0.0004089 0          0.000409 0           0.0004099 0          0.00041 1.5          0.0004109 1.5        0.000411 0           0.0004119 0          0.000412 0           0.0004129 0          0.000413 0           0.0004139 0          0.000414 1.5         0.0004149 1.5        0.000415 0           0.0004159 0          0.000416 0           0.0004169 0          0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.2          0.0005309 0.2        0.000531 0           0.0005319 0          0.000532 0.2         0.0005329 0.2        0.000533 0           0.0005339 0          0.000534 0.2         0.0005349 0.2        0.000535 0           0.0005359 0          0.000536 0.2         0.0005369 0.2        0.000537 0           0.0005379 0          0.000538 0.2         0.0005389 0.2        0.000539 0           0.0005399 0          0.00054 0.2          0.0005409 0.2        0.000541 0           0.0005419 0          0.000542 0.2         0.0005429 0.2        0.000543 0           0.0005439 0          0.000544 0.2         0.0005449 0.2        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_2 row_2_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.2          3.49e-05 0.2         3.5e-05 0            3.59e-05 0           3.6e-05 0.2          3.69e-05 0.2         3.7e-05 0            3.79e-05 0           3.8e-05 0.2          3.89e-05 0.2         3.9e-05 0            3.99e-05 0           4e-05 0.2            4.09e-05 0.2         4.1e-05 0            4.19e-05 0           4.2e-05 0.2          4.29e-05 0.2         4.3e-05 0            4.39e-05 0           4.4e-05 0.2          4.49e-05 0.2         4.5e-05 0            4.59e-05 0           4.6e-05 0.2          4.69e-05 0.2         4.7e-05 0            4.79e-05 0           4.8e-05 0.2          4.89e-05 0.2         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 1.5         0.0001629 1.5        0.000163 0           0.0001639 0          0.000164 0           0.0001649 0          0.000165 0           0.0001659 0          0.000166 1.5         0.0001669 1.5        0.000167 0           0.0001679 0          0.000168 0           0.0001689 0          0.000169 0           0.0001699 0          0.00017 1.5          0.0001709 1.5        0.000171 0           0.0001719 0          0.000172 0           0.0001729 0          0.000173 0           0.0001739 0          0.000174 1.5         0.0001749 1.5        0.000175 0           0.0001759 0          0.000176 0           0.0001769 0          0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.2          0.0002909 0.2        0.000291 0           0.0002919 0          0.000292 0.2         0.0002929 0.2        0.000293 0           0.0002939 0          0.000294 0.2         0.0002949 0.2        0.000295 0           0.0002959 0          0.000296 0.2         0.0002969 0.2        0.000297 0           0.0002979 0          0.000298 0.2         0.0002989 0.2        0.000299 0           0.0002999 0          0.0003 0.2           0.0003009 0.2        0.000301 0           0.0003019 0          0.000302 0.2         0.0003029 0.2        0.000303 0           0.0003039 0          0.000304 0.2         0.0003049 0.2        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0           0.0004189 0          0.000419 0           0.0004199 0          0.00042 1.5          0.0004209 1.5        0.000421 0           0.0004219 0          0.000422 0           0.0004229 0          0.000423 0           0.0004239 0          0.000424 1.5         0.0004249 1.5        0.000425 0           0.0004259 0          0.000426 0           0.0004269 0          0.000427 0           0.0004279 0          0.000428 1.5         0.0004289 1.5        0.000429 0           0.0004299 0          0.00043 0            0.0004309 0          0.000431 0           0.0004319 0          0.000432 1.5         0.0004329 1.5        0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.2         0.0005469 0.2        0.000547 0           0.0005479 0          0.000548 0.2         0.0005489 0.2        0.000549 0           0.0005499 0          0.00055 0.2          0.0005509 0.2        0.000551 0           0.0005519 0          0.000552 0.2         0.0005529 0.2        0.000553 0           0.0005539 0          0.000554 0.2         0.0005549 0.2        0.000555 0           0.0005559 0          0.000556 0.2         0.0005569 0.2        0.000557 0           0.0005579 0          0.000558 0.2         0.0005589 0.2        0.000559 0           0.0005599 0          0.00056 0.2          0.0005609 0.2        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_3 row_3_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.2            5.09e-05 0.2         5.1e-05 0            5.19e-05 0           5.2e-05 0.2          5.29e-05 0.2         5.3e-05 0            5.39e-05 0           5.4e-05 0.2          5.49e-05 0.2         5.5e-05 0            5.59e-05 0           5.6e-05 0.2          5.69e-05 0.2         5.7e-05 0            5.79e-05 0           5.8e-05 0.2          5.89e-05 0.2         5.9e-05 0            5.99e-05 0           6e-05 0.2            6.09e-05 0.2         6.1e-05 0            6.19e-05 0           6.2e-05 0.2          6.29e-05 0.2         6.3e-05 0            6.39e-05 0           6.4e-05 0.2          6.49e-05 0.2         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0           0.0001789 0          0.000179 0           0.0001799 0          0.00018 1.5          0.0001809 1.5        0.000181 0           0.0001819 0          0.000182 0           0.0001829 0          0.000183 0           0.0001839 0          0.000184 1.5         0.0001849 1.5        0.000185 0           0.0001859 0          0.000186 0           0.0001869 0          0.000187 0           0.0001879 0          0.000188 1.5         0.0001889 1.5        0.000189 0           0.0001899 0          0.00019 0            0.0001909 0          0.000191 0           0.0001919 0          0.000192 1.5         0.0001929 1.5        0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.2         0.0003069 0.2        0.000307 0           0.0003079 0          0.000308 0.2         0.0003089 0.2        0.000309 0           0.0003099 0          0.00031 0.2          0.0003109 0.2        0.000311 0           0.0003119 0          0.000312 0.2         0.0003129 0.2        0.000313 0           0.0003139 0          0.000314 0.2         0.0003149 0.2        0.000315 0           0.0003159 0          0.000316 0.2         0.0003169 0.2        0.000317 0           0.0003179 0          0.000318 0.2         0.0003189 0.2        0.000319 0           0.0003199 0          0.00032 0.2          0.0003209 0.2        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 1.5         0.0004349 1.5        0.000435 0           0.0004359 0          0.000436 0           0.0004369 0          0.000437 0           0.0004379 0          0.000438 1.5         0.0004389 1.5        0.000439 0           0.0004399 0          0.00044 0            0.0004409 0          0.000441 0           0.0004419 0          0.000442 1.5         0.0004429 1.5        0.000443 0           0.0004439 0          0.000444 0           0.0004449 0          0.000445 0           0.0004459 0          0.000446 1.5         0.0004469 1.5        0.000447 0           0.0004479 0          0.000448 0           0.0004489 0          0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.2         0.0005629 0.2        0.000563 0           0.0005639 0          0.000564 0.2         0.0005649 0.2        0.000565 0           0.0005659 0          0.000566 0.2         0.0005669 0.2        0.000567 0           0.0005679 0          0.000568 0.2         0.0005689 0.2        0.000569 0           0.0005699 0          0.00057 0.2          0.0005709 0.2        0.000571 0           0.0005719 0          0.000572 0.2         0.0005729 0.2        0.000573 0           0.0005739 0          0.000574 0.2         0.0005749 0.2        0.000575 0           0.0005759 0          0.000576 0.2         0.0005769 0.2        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_4 row_4_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.2          6.69e-05 0.2         6.7e-05 0            6.79e-05 0           6.8e-05 0.2          6.89e-05 0.2         6.9e-05 0            6.99e-05 0           7e-05 0.2            7.09e-05 0.2         7.1e-05 0            7.19e-05 0           7.2e-05 0.2          7.29e-05 0.2         7.3e-05 0            7.39e-05 0           7.4e-05 0.2          7.49e-05 0.2         7.5e-05 0            7.59e-05 0           7.6e-05 0.2          7.69e-05 0.2         7.7e-05 0            7.79e-05 0           7.8e-05 0.2          7.89e-05 0.2         7.9e-05 0            7.99e-05 0           8e-05 0.2            8.09e-05 0.2         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 1.5         0.0001949 1.5        0.000195 0           0.0001959 0          0.000196 0           0.0001969 0          0.000197 0           0.0001979 0          0.000198 1.5         0.0001989 1.5        0.000199 0           0.0001999 0          0.0002 0             0.0002009 0          0.000201 0           0.0002019 0          0.000202 1.5         0.0002029 1.5        0.000203 0           0.0002039 0          0.000204 0           0.0002049 0          0.000205 0           0.0002059 0          0.000206 1.5         0.0002069 1.5        0.000207 0           0.0002079 0          0.000208 0           0.0002089 0          0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.2         0.0003229 0.2        0.000323 0           0.0003239 0          0.000324 0.2         0.0003249 0.2        0.000325 0           0.0003259 0          0.000326 0.2         0.0003269 0.2        0.000327 0           0.0003279 0          0.000328 0.2         0.0003289 0.2        0.000329 0           0.0003299 0          0.00033 0.2          0.0003309 0.2        0.000331 0           0.0003319 0          0.000332 0.2         0.0003329 0.2        0.000333 0           0.0003339 0          0.000334 0.2         0.0003349 0.2        0.000335 0           0.0003359 0          0.000336 0.2         0.0003369 0.2        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0            0.0004509 0          0.000451 0           0.0004519 0          0.000452 1.5         0.0004529 1.5        0.000453 0           0.0004539 0          0.000454 0           0.0004549 0          0.000455 0           0.0004559 0          0.000456 1.5         0.0004569 1.5        0.000457 0           0.0004579 0          0.000458 0           0.0004589 0          0.000459 0           0.0004599 0          0.00046 1.5          0.0004609 1.5        0.000461 0           0.0004619 0          0.000462 0           0.0004629 0          0.000463 0           0.0004639 0          0.000464 1.5         0.0004649 1.5        0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.2         0.0005789 0.2        0.000579 0           0.0005799 0          0.00058 0.2          0.0005809 0.2        0.000581 0           0.0005819 0          0.000582 0.2         0.0005829 0.2        0.000583 0           0.0005839 0          0.000584 0.2         0.0005849 0.2        0.000585 0           0.0005859 0          0.000586 0.2         0.0005869 0.2        0.000587 0           0.0005879 0          0.000588 0.2         0.0005889 0.2        0.000589 0           0.0005899 0          0.00059 0.2          0.0005909 0.2        0.000591 0           0.0005919 0          0.000592 0.2         0.0005929 0.2        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_5 row_5_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.2          8.29e-05 0.2         8.3e-05 0            8.39e-05 0           8.4e-05 0.2          8.49e-05 0.2         8.5e-05 0            8.59e-05 0           8.6e-05 0.2          8.69e-05 0.2         8.7e-05 0            8.79e-05 0           8.8e-05 0.2          8.89e-05 0.2         8.9e-05 0            8.99e-05 0           9e-05 0.2            9.09e-05 0.2         9.1e-05 0            9.19e-05 0           9.2e-05 0.2          9.29e-05 0.2         9.3e-05 0            9.39e-05 0           9.4e-05 0.2          9.49e-05 0.2         9.5e-05 0            9.59e-05 0           9.6e-05 0.2          9.69e-05 0.2         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0            0.0002109 0          0.000211 0           0.0002119 0          0.000212 1.5         0.0002129 1.5        0.000213 0           0.0002139 0          0.000214 0           0.0002149 0          0.000215 0           0.0002159 0          0.000216 1.5         0.0002169 1.5        0.000217 0           0.0002179 0          0.000218 0           0.0002189 0          0.000219 0           0.0002199 0          0.00022 1.5          0.0002209 1.5        0.000221 0           0.0002219 0          0.000222 0           0.0002229 0          0.000223 0           0.0002239 0          0.000224 1.5         0.0002249 1.5        0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.2         0.0003389 0.2        0.000339 0           0.0003399 0          0.00034 0.2          0.0003409 0.2        0.000341 0           0.0003419 0          0.000342 0.2         0.0003429 0.2        0.000343 0           0.0003439 0          0.000344 0.2         0.0003449 0.2        0.000345 0           0.0003459 0          0.000346 0.2         0.0003469 0.2        0.000347 0           0.0003479 0          0.000348 0.2         0.0003489 0.2        0.000349 0           0.0003499 0          0.00035 0.2          0.0003509 0.2        0.000351 0           0.0003519 0          0.000352 0.2         0.0003529 0.2        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 1.5         0.0004669 1.5        0.000467 0           0.0004679 0          0.000468 0           0.0004689 0          0.000469 0           0.0004699 0          0.00047 1.5          0.0004709 1.5        0.000471 0           0.0004719 0          0.000472 0           0.0004729 0          0.000473 0           0.0004739 0          0.000474 1.5         0.0004749 1.5        0.000475 0           0.0004759 0          0.000476 0           0.0004769 0          0.000477 0           0.0004779 0          0.000478 1.5         0.0004789 1.5        0.000479 0           0.0004799 0          0.00048 0            0.0004809 0          0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.2         0.0005949 0.2        0.000595 0           0.0005959 0          0.000596 0.2         0.0005969 0.2        0.000597 0           0.0005979 0          0.000598 0.2         0.0005989 0.2        0.000599 0           0.0005999 0          0.0006 0.2           0.0006009 0.2        0.000601 0           0.0006019 0          0.000602 0.2         0.0006029 0.2        0.000603 0           0.0006039 0          0.000604 0.2         0.0006049 0.2        0.000605 0           0.0006059 0          0.000606 0.2         0.0006069 0.2        0.000607 0           0.0006079 0          0.000608 0.2         0.0006089 0.2        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_6 row_6_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.2          9.89e-05 0.2         9.9e-05 0            9.99e-05 0           0.0001 0.2           0.0001009 0.2        0.000101 0           0.0001019 0          0.000102 0.2         0.0001029 0.2        0.000103 0           0.0001039 0          0.000104 0.2         0.0001049 0.2        0.000105 0           0.0001059 0          0.000106 0.2         0.0001069 0.2        0.000107 0           0.0001079 0          0.000108 0.2         0.0001089 0.2        0.000109 0           0.0001099 0          0.00011 0.2          0.0001109 0.2        0.000111 0           0.0001119 0          0.000112 0.2         0.0001129 0.2        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 1.5         0.0002269 1.5        0.000227 0           0.0002279 0          0.000228 0           0.0002289 0          0.000229 0           0.0002299 0          0.00023 1.5          0.0002309 1.5        0.000231 0           0.0002319 0          0.000232 0           0.0002329 0          0.000233 0           0.0002339 0          0.000234 1.5         0.0002349 1.5        0.000235 0           0.0002359 0          0.000236 0           0.0002369 0          0.000237 0           0.0002379 0          0.000238 1.5         0.0002389 1.5        0.000239 0           0.0002399 0          0.00024 0            0.0002409 0          0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.2         0.0003549 0.2        0.000355 0           0.0003559 0          0.000356 0.2         0.0003569 0.2        0.000357 0           0.0003579 0          0.000358 0.2         0.0003589 0.2        0.000359 0           0.0003599 0          0.00036 0.2          0.0003609 0.2        0.000361 0           0.0003619 0          0.000362 0.2         0.0003629 0.2        0.000363 0           0.0003639 0          0.000364 0.2         0.0003649 0.2        0.000365 0           0.0003659 0          0.000366 0.2         0.0003669 0.2        0.000367 0           0.0003679 0          0.000368 0.2         0.0003689 0.2        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0           0.0004829 0          0.000483 0           0.0004839 0          0.000484 1.5         0.0004849 1.5        0.000485 0           0.0004859 0          0.000486 0           0.0004869 0          0.000487 0           0.0004879 0          0.000488 1.5         0.0004889 1.5        0.000489 0           0.0004899 0          0.00049 0            0.0004909 0          0.000491 0           0.0004919 0          0.000492 1.5         0.0004929 1.5        0.000493 0           0.0004939 0          0.000494 0           0.0004949 0          0.000495 0           0.0004959 0          0.000496 1.5         0.0004969 1.5        0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.2          0.0006109 0.2        0.000611 0           0.0006119 0          0.000612 0.2         0.0006129 0.2        0.000613 0           0.0006139 0          0.000614 0.2         0.0006149 0.2        0.000615 0           0.0006159 0          0.000616 0.2         0.0006169 0.2        0.000617 0           0.0006179 0          0.000618 0.2         0.0006189 0.2        0.000619 0           0.0006199 0          0.00062 0.2          0.0006209 0.2        0.000621 0           0.0006219 0          0.000622 0.2         0.0006229 0.2        0.000623 0           0.0006239 0          0.000624 0.2         0.0006249 0.2        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vrow_7 row_7_0 0 PWLZ(0 0                  9e-07 0              1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.2         0.0001149 0.2        0.000115 0           0.0001159 0          0.000116 0.2         0.0001169 0.2        0.000117 0           0.0001179 0          0.000118 0.2         0.0001189 0.2        0.000119 0           0.0001199 0          0.00012 0.2          0.0001209 0.2        0.000121 0           0.0001219 0          0.000122 0.2         0.0001229 0.2        0.000123 0           0.0001239 0          0.000124 0.2         0.0001249 0.2        0.000125 0           0.0001259 0          0.000126 0.2         0.0001269 0.2        0.000127 0           0.0001279 0          0.000128 0.2         0.0001289 0.2        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0           0.0002429 0          0.000243 0           0.0002439 0          0.000244 1.5         0.0002449 1.5        0.000245 0           0.0002459 0          0.000246 0           0.0002469 0          0.000247 0           0.0002479 0          0.000248 1.5         0.0002489 1.5        0.000249 0           0.0002499 0          0.00025 0            0.0002509 0          0.000251 0           0.0002519 0          0.000252 1.5         0.0002529 1.5        0.000253 0           0.0002539 0          0.000254 0           0.0002549 0          0.000255 0           0.0002559 0          0.000256 1.5         0.0002569 1.5        0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.2          0.0003709 0.2        0.000371 0           0.0003719 0          0.000372 0.2         0.0003729 0.2        0.000373 0           0.0003739 0          0.000374 0.2         0.0003749 0.2        0.000375 0           0.0003759 0          0.000376 0.2         0.0003769 0.2        0.000377 0           0.0003779 0          0.000378 0.2         0.0003789 0.2        0.000379 0           0.0003799 0          0.00038 0.2          0.0003809 0.2        0.000381 0           0.0003819 0          0.000382 0.2         0.0003829 0.2        0.000383 0           0.0003839 0          0.000384 0.2         0.0003849 0.2        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 1.5         0.0004989 1.5        0.000499 0           0.0004999 0          0.0005 0             0.0005009 0          0.000501 0           0.0005019 0          0.000502 1.5         0.0005029 1.5        0.000503 0           0.0005039 0          0.000504 0           0.0005049 0          0.000505 0           0.0005059 0          0.000506 1.5         0.0005069 1.5        0.000507 0           0.0005079 0          0.000508 0           0.0005089 0          0.000509 0           0.0005099 0          0.00051 1.5          0.0005109 1.5        0.000511 0           0.0005119 0          0.000512 0           0.0005129 0          0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.2         0.0006269 0.2        0.000627 0           0.0006279 0          0.000628 0.2         0.0006289 0.2        0.000629 0           0.0006299 0          0.00063 0.2          0.0006309 0.2        0.000631 0           0.0006319 0          0.000632 0.2         0.0006329 0.2        0.000633 0           0.0006339 0          0.000634 0.2         0.0006349 0.2        0.000635 0           0.0006359 0          0.000636 0.2         0.0006369 0.2        0.000637 0           0.0006379 0          0.000638 0.2         0.0006389 0.2        0.000639 0           0.0006399 0          0.00064 0.2          0.0006409 0.2        0.000641 0           0.0006419 0         )
Vcol_0 col_0_0 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0              2.9e-06 0            3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0            1.89e-05 0           1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0            3.49e-05 0           3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0              5.09e-05 0           5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0            6.69e-05 0           6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0            8.29e-05 0           8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0            9.89e-05 0           9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0           0.0001149 0          0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0            0.0001309 0          0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 1.5         0.0001469 1.5        0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0           0.0001629 0          0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 1.5         0.0001789 1.5        0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0           0.0001949 0          0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 1.5          0.0002109 1.5        0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0           0.0002269 0          0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 1.5         0.0002429 1.5        0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0           0.0002589 0          0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0           0.0002749 0          0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0            0.0002909 0          0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0           0.0003069 0          0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0           0.0003229 0          0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0           0.0003389 0          0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0           0.0003549 0          0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0            0.0003709 0          0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 1.5         0.0003869 1.5        0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0           0.0004029 0          0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 1.5         0.0004189 1.5        0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0           0.0004349 0          0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 1.5          0.0004509 1.5        0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0           0.0004669 0          0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 1.5         0.0004829 1.5        0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0           0.0004989 0          0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0           0.0005149 0          0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0            0.0005309 0          0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0           0.0005469 0          0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0           0.0005629 0          0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0           0.0005789 0          0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0           0.0005949 0          0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0            0.0006109 0          0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0           0.0006269 0          0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_1 col_0_1 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0              4.9e-06 0            5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0              2.09e-05 0           2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0            3.69e-05 0           3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0            5.29e-05 0           5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0            6.89e-05 0           6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0            8.49e-05 0           8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0             0.0001009 0          0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0           0.0001169 0          0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 1.5         0.0001329 1.5        0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0           0.0001489 0          0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 1.5         0.0001649 1.5        0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0            0.0001809 0          0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 1.5         0.0001969 1.5        0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0           0.0002129 0          0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 1.5         0.0002289 1.5        0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0           0.0002449 0          0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0            0.0002609 0          0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0           0.0002769 0          0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0           0.0002929 0          0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0           0.0003089 0          0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0           0.0003249 0          0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0            0.0003409 0          0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0           0.0003569 0          0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0           0.0003729 0          0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0           0.0003889 0          0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 1.5         0.0004049 1.5        0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0            0.0004209 0          0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 1.5         0.0004369 1.5        0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0           0.0004529 0          0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 1.5         0.0004689 1.5        0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0           0.0004849 0          0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 1.5           0.0005009 1.5        0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0           0.0005169 0          0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0           0.0005329 0          0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0           0.0005489 0          0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0           0.0005649 0          0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0            0.0005809 0          0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0           0.0005969 0          0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0           0.0006129 0          0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0           0.0006289 0          0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_2 col_0_2 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0              6.9e-06 0            7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0            2.29e-05 0           2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0            3.89e-05 0           3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0            5.49e-05 0           5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0              7.09e-05 0           7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0            8.69e-05 0           8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0           0.0001029 0          0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0           0.0001189 0          0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0           0.0001349 0          0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 1.5          0.0001509 1.5        0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0           0.0001669 0          0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 1.5         0.0001829 1.5        0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0           0.0001989 0          0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 1.5         0.0002149 1.5        0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0            0.0002309 0          0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 1.5         0.0002469 1.5        0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0           0.0002629 0          0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0           0.0002789 0          0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0           0.0002949 0          0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0            0.0003109 0          0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0           0.0003269 0          0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0           0.0003429 0          0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0           0.0003589 0          0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0           0.0003749 0          0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 1.5          0.0003909 1.5        0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0           0.0004069 0          0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 1.5         0.0004229 1.5        0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0           0.0004389 0          0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 1.5         0.0004549 1.5        0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0            0.0004709 0          0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 1.5         0.0004869 1.5        0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0           0.0005029 0          0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0           0.0005189 0          0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0           0.0005349 0          0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0            0.0005509 0          0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0           0.0005669 0          0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0           0.0005829 0          0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0           0.0005989 0          0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0           0.0006149 0          0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0            0.0006309 0          0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_3 col_0_3 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0              8.9e-06 0            9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0            2.49e-05 0           2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0              4.09e-05 0           4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0            5.69e-05 0           5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0            7.29e-05 0           7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0            8.89e-05 0           8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0           0.0001049 0          0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0            0.0001209 0          0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 1.5         0.0001369 1.5        0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0           0.0001529 0          0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 1.5         0.0001689 1.5        0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0           0.0001849 0          0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 1.5           0.0002009 1.5        0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0           0.0002169 0          0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 1.5         0.0002329 1.5        0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0           0.0002489 0          0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0           0.0002649 0          0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0            0.0002809 0          0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0           0.0002969 0          0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0           0.0003129 0          0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0           0.0003289 0          0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0           0.0003449 0          0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0            0.0003609 0          0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0           0.0003769 0          0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0           0.0003929 0          0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 1.5         0.0004089 1.5        0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0           0.0004249 0          0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 1.5          0.0004409 1.5        0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0           0.0004569 0          0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 1.5         0.0004729 1.5        0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0           0.0004889 0          0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 1.5         0.0005049 1.5        0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0            0.0005209 0          0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0           0.0005369 0          0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0           0.0005529 0          0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0           0.0005689 0          0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0           0.0005849 0          0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0             0.0006009 0          0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0           0.0006169 0          0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0           0.0006329 0          0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_4 col_0_4 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0              1.09e-05 0           1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0            2.69e-05 0           2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0            4.29e-05 0           4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0            5.89e-05 0           5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0            7.49e-05 0           7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0              9.09e-05 0           9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0           0.0001069 0          0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0           0.0001229 0          0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0           0.0001389 0          0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 1.5         0.0001549 1.5        0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0            0.0001709 0          0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 1.5         0.0001869 1.5        0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0           0.0002029 0          0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 1.5         0.0002189 1.5        0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0           0.0002349 0          0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 1.5          0.0002509 1.5        0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0           0.0002669 0          0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0           0.0002829 0          0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0           0.0002989 0          0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0           0.0003149 0          0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0            0.0003309 0          0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0           0.0003469 0          0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0           0.0003629 0          0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0           0.0003789 0          0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 1.5         0.0003949 1.5        0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0            0.0004109 0          0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 1.5         0.0004269 1.5        0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0           0.0004429 0          0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 1.5         0.0004589 1.5        0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0           0.0004749 0          0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 1.5          0.0004909 1.5        0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0           0.0005069 0          0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0           0.0005229 0          0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0           0.0005389 0          0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0           0.0005549 0          0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0            0.0005709 0          0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0           0.0005869 0          0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0           0.0006029 0          0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0           0.0006189 0          0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0           0.0006349 0          0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_5 col_0_5 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0            1.29e-05 0           1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0            2.89e-05 0           2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0            4.49e-05 0           4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0              6.09e-05 0           6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0            7.69e-05 0           7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0            9.29e-05 0           9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0           0.0001089 0          0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0           0.0001249 0          0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 1.5          0.0001409 1.5        0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0           0.0001569 0          0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 1.5         0.0001729 1.5        0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0           0.0001889 0          0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 1.5         0.0002049 1.5        0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0            0.0002209 0          0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 1.5         0.0002369 1.5        0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0           0.0002529 0          0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0           0.0002689 0          0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0           0.0002849 0          0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0             0.0003009 0          0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0           0.0003169 0          0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0           0.0003329 0          0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0           0.0003489 0          0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0           0.0003649 0          0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0            0.0003809 0          0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0           0.0003969 0          0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 1.5         0.0004129 1.5        0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0           0.0004289 0          0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 1.5         0.0004449 1.5        0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0            0.0004609 0          0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 1.5         0.0004769 1.5        0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0           0.0004929 0          0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 1.5         0.0005089 1.5        0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0           0.0005249 0          0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0            0.0005409 0          0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0           0.0005569 0          0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0           0.0005729 0          0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0           0.0005889 0          0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0           0.0006049 0          0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0            0.0006209 0          0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0           0.0006369 0          0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_6 col_0_6 0 PWLZ(0 0.0                9e-07 0.0            1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0            1.49e-05 0           1.5e-05 0            1.59e-05 0           1.6e-05 0.1          1.69e-05 0.1         1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0              3.09e-05 0           3.1e-05 0            3.19e-05 0           3.2e-05 0.1          3.29e-05 0.1         3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0            4.69e-05 0           4.7e-05 0            4.79e-05 0           4.8e-05 0.1          4.89e-05 0.1         4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0            6.29e-05 0           6.3e-05 0            6.39e-05 0           6.4e-05 0.1          6.49e-05 0.1         6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0            7.89e-05 0           7.9e-05 0            7.99e-05 0           8e-05 0.1            8.09e-05 0.1         8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0            9.49e-05 0           9.5e-05 0            9.59e-05 0           9.6e-05 0.1          9.69e-05 0.1         9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0            0.0001109 0          0.000111 0           0.0001119 0          0.000112 0.1         0.0001129 0.1        0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0           0.0001269 0          0.000127 0           0.0001279 0          0.000128 0.1         0.0001289 0.1        0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0           0.0001429 0          0.000143 0           0.0001439 0          0.000144 0.75        0.0001449 0.75       0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 1.5         0.0001589 1.5        0.000159 0           0.0001599 0          0.00016 0.75         0.0001609 0.75       0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0           0.0001749 0          0.000175 0           0.0001759 0          0.000176 0.75        0.0001769 0.75       0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 1.5          0.0001909 1.5        0.000191 0           0.0001919 0          0.000192 0.75        0.0001929 0.75       0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0           0.0002069 0          0.000207 0           0.0002079 0          0.000208 0.75        0.0002089 0.75       0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 1.5         0.0002229 1.5        0.000223 0           0.0002239 0          0.000224 0.75        0.0002249 0.75       0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0           0.0002389 0          0.000239 0           0.0002399 0          0.00024 0.75         0.0002409 0.75       0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 1.5         0.0002549 1.5        0.000255 0           0.0002559 0          0.000256 0.75        0.0002569 0.75       0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0            0.0002709 0          0.000271 0           0.0002719 0          0.000272 0.1         0.0002729 0.1        0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0           0.0002869 0          0.000287 0           0.0002879 0          0.000288 0.1         0.0002889 0.1        0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0           0.0003029 0          0.000303 0           0.0003039 0          0.000304 0.1         0.0003049 0.1        0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0           0.0003189 0          0.000319 0           0.0003199 0          0.00032 0.1          0.0003209 0.1        0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0           0.0003349 0          0.000335 0           0.0003359 0          0.000336 0.1         0.0003369 0.1        0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0            0.0003509 0          0.000351 0           0.0003519 0          0.000352 0.1         0.0003529 0.1        0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0           0.0003669 0          0.000367 0           0.0003679 0          0.000368 0.1         0.0003689 0.1        0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0           0.0003829 0          0.000383 0           0.0003839 0          0.000384 0.1         0.0003849 0.1        0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 1.5         0.0003989 1.5        0.000399 0           0.0003999 0          0.0004 0.75          0.0004009 0.75       0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0           0.0004149 0          0.000415 0           0.0004159 0          0.000416 0.75        0.0004169 0.75       0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 1.5          0.0004309 1.5        0.000431 0           0.0004319 0          0.000432 0.75        0.0004329 0.75       0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0           0.0004469 0          0.000447 0           0.0004479 0          0.000448 0.75        0.0004489 0.75       0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 1.5         0.0004629 1.5        0.000463 0           0.0004639 0          0.000464 0.75        0.0004649 0.75       0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0           0.0004789 0          0.000479 0           0.0004799 0          0.00048 0.75         0.0004809 0.75       0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 1.5         0.0004949 1.5        0.000495 0           0.0004959 0          0.000496 0.75        0.0004969 0.75       0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0            0.0005109 0          0.000511 0           0.0005119 0          0.000512 0.75        0.0005129 0.75       0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0           0.0005269 0          0.000527 0           0.0005279 0          0.000528 0.1         0.0005289 0.1        0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0           0.0005429 0          0.000543 0           0.0005439 0          0.000544 0.1         0.0005449 0.1        0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0           0.0005589 0          0.000559 0           0.0005599 0          0.00056 0.1          0.0005609 0.1        0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0           0.0005749 0          0.000575 0           0.0005759 0          0.000576 0.1         0.0005769 0.1        0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0            0.0005909 0          0.000591 0           0.0005919 0          0.000592 0.1         0.0005929 0.1        0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0           0.0006069 0          0.000607 0           0.0006079 0          0.000608 0.1         0.0006089 0.1        0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0           0.0006229 0          0.000623 0           0.0006239 0          0.000624 0.1         0.0006249 0.1        0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0           0.0006389 0          0.000639 0           0.0006399 0          0.00064 0.1          0.0006409 0.1        0.000641 0           0.0006419 0         )
Vcol_7 col_0_7 0 PWLZ(0 0                  9e-07 0              1e-06 0              1.9e-06 0            2e-06 0.1            2.9e-06 0.1          3e-06 0              3.9e-06 0            4e-06 0.1            4.9e-06 0.1          5e-06 0              5.9e-06 0            6e-06 0.1            6.9e-06 0.1          7e-06 0              7.9e-06 0            8e-06 0.1            8.9e-06 0.1          9e-06 0              9.9e-06 0            1e-05 0.1            1.09e-05 0.1         1.1e-05 0            1.19e-05 0           1.2e-05 0.1          1.29e-05 0.1         1.3e-05 0            1.39e-05 0           1.4e-05 0.1          1.49e-05 0.1         1.5e-05 0            1.59e-05 0           1.6e-05 0            1.69e-05 0           1.7e-05 0            1.79e-05 0           1.8e-05 0.1          1.89e-05 0.1         1.9e-05 0            1.99e-05 0           2e-05 0.1            2.09e-05 0.1         2.1e-05 0            2.19e-05 0           2.2e-05 0.1          2.29e-05 0.1         2.3e-05 0            2.39e-05 0           2.4e-05 0.1          2.49e-05 0.1         2.5e-05 0            2.59e-05 0           2.6e-05 0.1          2.69e-05 0.1         2.7e-05 0            2.79e-05 0           2.8e-05 0.1          2.89e-05 0.1         2.9e-05 0            2.99e-05 0           3e-05 0.1            3.09e-05 0.1         3.1e-05 0            3.19e-05 0           3.2e-05 0            3.29e-05 0           3.3e-05 0            3.39e-05 0           3.4e-05 0.1          3.49e-05 0.1         3.5e-05 0            3.59e-05 0           3.6e-05 0.1          3.69e-05 0.1         3.7e-05 0            3.79e-05 0           3.8e-05 0.1          3.89e-05 0.1         3.9e-05 0            3.99e-05 0           4e-05 0.1            4.09e-05 0.1         4.1e-05 0            4.19e-05 0           4.2e-05 0.1          4.29e-05 0.1         4.3e-05 0            4.39e-05 0           4.4e-05 0.1          4.49e-05 0.1         4.5e-05 0            4.59e-05 0           4.6e-05 0.1          4.69e-05 0.1         4.7e-05 0            4.79e-05 0           4.8e-05 0            4.89e-05 0           4.9e-05 0            4.99e-05 0           5e-05 0.1            5.09e-05 0.1         5.1e-05 0            5.19e-05 0           5.2e-05 0.1          5.29e-05 0.1         5.3e-05 0            5.39e-05 0           5.4e-05 0.1          5.49e-05 0.1         5.5e-05 0            5.59e-05 0           5.6e-05 0.1          5.69e-05 0.1         5.7e-05 0            5.79e-05 0           5.8e-05 0.1          5.89e-05 0.1         5.9e-05 0            5.99e-05 0           6e-05 0.1            6.09e-05 0.1         6.1e-05 0            6.19e-05 0           6.2e-05 0.1          6.29e-05 0.1         6.3e-05 0            6.39e-05 0           6.4e-05 0            6.49e-05 0           6.5e-05 0            6.59e-05 0           6.6e-05 0.1          6.69e-05 0.1         6.7e-05 0            6.79e-05 0           6.8e-05 0.1          6.89e-05 0.1         6.9e-05 0            6.99e-05 0           7e-05 0.1            7.09e-05 0.1         7.1e-05 0            7.19e-05 0           7.2e-05 0.1          7.29e-05 0.1         7.3e-05 0            7.39e-05 0           7.4e-05 0.1          7.49e-05 0.1         7.5e-05 0            7.59e-05 0           7.6e-05 0.1          7.69e-05 0.1         7.7e-05 0            7.79e-05 0           7.8e-05 0.1          7.89e-05 0.1         7.9e-05 0            7.99e-05 0           8e-05 0              8.09e-05 0           8.1e-05 0            8.19e-05 0           8.2e-05 0.1          8.29e-05 0.1         8.3e-05 0            8.39e-05 0           8.4e-05 0.1          8.49e-05 0.1         8.5e-05 0            8.59e-05 0           8.6e-05 0.1          8.69e-05 0.1         8.7e-05 0            8.79e-05 0           8.8e-05 0.1          8.89e-05 0.1         8.9e-05 0            8.99e-05 0           9e-05 0.1            9.09e-05 0.1         9.1e-05 0            9.19e-05 0           9.2e-05 0.1          9.29e-05 0.1         9.3e-05 0            9.39e-05 0           9.4e-05 0.1          9.49e-05 0.1         9.5e-05 0            9.59e-05 0           9.6e-05 0            9.69e-05 0           9.7e-05 0            9.79e-05 0           9.8e-05 0.1          9.89e-05 0.1         9.9e-05 0            9.99e-05 0           0.0001 0.1           0.0001009 0.1        0.000101 0           0.0001019 0          0.000102 0.1         0.0001029 0.1        0.000103 0           0.0001039 0          0.000104 0.1         0.0001049 0.1        0.000105 0           0.0001059 0          0.000106 0.1         0.0001069 0.1        0.000107 0           0.0001079 0          0.000108 0.1         0.0001089 0.1        0.000109 0           0.0001099 0          0.00011 0.1          0.0001109 0.1        0.000111 0           0.0001119 0          0.000112 0           0.0001129 0          0.000113 0           0.0001139 0          0.000114 0.1         0.0001149 0.1        0.000115 0           0.0001159 0          0.000116 0.1         0.0001169 0.1        0.000117 0           0.0001179 0          0.000118 0.1         0.0001189 0.1        0.000119 0           0.0001199 0          0.00012 0.1          0.0001209 0.1        0.000121 0           0.0001219 0          0.000122 0.1         0.0001229 0.1        0.000123 0           0.0001239 0          0.000124 0.1         0.0001249 0.1        0.000125 0           0.0001259 0          0.000126 0.1         0.0001269 0.1        0.000127 0           0.0001279 0          0.000128 0           0.0001289 0          0.000129 0           0.0001299 0          0.00013 0.75         0.0001309 0.75       0.000131 0           0.0001319 0          0.000132 0.75        0.0001329 0.75       0.000133 0           0.0001339 0          0.000134 0.75        0.0001349 0.75       0.000135 0           0.0001359 0          0.000136 0.75        0.0001369 0.75       0.000137 0           0.0001379 0          0.000138 0.75        0.0001389 0.75       0.000139 0           0.0001399 0          0.00014 0.75         0.0001409 0.75       0.000141 0           0.0001419 0          0.000142 0.75        0.0001429 0.75       0.000143 0           0.0001439 0          0.000144 1.5         0.0001449 1.5        0.000145 0           0.0001459 0          0.000146 0.75        0.0001469 0.75       0.000147 0           0.0001479 0          0.000148 0.75        0.0001489 0.75       0.000149 0           0.0001499 0          0.00015 0.75         0.0001509 0.75       0.000151 0           0.0001519 0          0.000152 0.75        0.0001529 0.75       0.000153 0           0.0001539 0          0.000154 0.75        0.0001549 0.75       0.000155 0           0.0001559 0          0.000156 0.75        0.0001569 0.75       0.000157 0           0.0001579 0          0.000158 0.75        0.0001589 0.75       0.000159 0           0.0001599 0          0.00016 0            0.0001609 0          0.000161 0           0.0001619 0          0.000162 0.75        0.0001629 0.75       0.000163 0           0.0001639 0          0.000164 0.75        0.0001649 0.75       0.000165 0           0.0001659 0          0.000166 0.75        0.0001669 0.75       0.000167 0           0.0001679 0          0.000168 0.75        0.0001689 0.75       0.000169 0           0.0001699 0          0.00017 0.75         0.0001709 0.75       0.000171 0           0.0001719 0          0.000172 0.75        0.0001729 0.75       0.000173 0           0.0001739 0          0.000174 0.75        0.0001749 0.75       0.000175 0           0.0001759 0          0.000176 1.5         0.0001769 1.5        0.000177 0           0.0001779 0          0.000178 0.75        0.0001789 0.75       0.000179 0           0.0001799 0          0.00018 0.75         0.0001809 0.75       0.000181 0           0.0001819 0          0.000182 0.75        0.0001829 0.75       0.000183 0           0.0001839 0          0.000184 0.75        0.0001849 0.75       0.000185 0           0.0001859 0          0.000186 0.75        0.0001869 0.75       0.000187 0           0.0001879 0          0.000188 0.75        0.0001889 0.75       0.000189 0           0.0001899 0          0.00019 0.75         0.0001909 0.75       0.000191 0           0.0001919 0          0.000192 0           0.0001929 0          0.000193 0           0.0001939 0          0.000194 0.75        0.0001949 0.75       0.000195 0           0.0001959 0          0.000196 0.75        0.0001969 0.75       0.000197 0           0.0001979 0          0.000198 0.75        0.0001989 0.75       0.000199 0           0.0001999 0          0.0002 0.75          0.0002009 0.75       0.000201 0           0.0002019 0          0.000202 0.75        0.0002029 0.75       0.000203 0           0.0002039 0          0.000204 0.75        0.0002049 0.75       0.000205 0           0.0002059 0          0.000206 0.75        0.0002069 0.75       0.000207 0           0.0002079 0          0.000208 1.5         0.0002089 1.5        0.000209 0           0.0002099 0          0.00021 0.75         0.0002109 0.75       0.000211 0           0.0002119 0          0.000212 0.75        0.0002129 0.75       0.000213 0           0.0002139 0          0.000214 0.75        0.0002149 0.75       0.000215 0           0.0002159 0          0.000216 0.75        0.0002169 0.75       0.000217 0           0.0002179 0          0.000218 0.75        0.0002189 0.75       0.000219 0           0.0002199 0          0.00022 0.75         0.0002209 0.75       0.000221 0           0.0002219 0          0.000222 0.75        0.0002229 0.75       0.000223 0           0.0002239 0          0.000224 0           0.0002249 0          0.000225 0           0.0002259 0          0.000226 0.75        0.0002269 0.75       0.000227 0           0.0002279 0          0.000228 0.75        0.0002289 0.75       0.000229 0           0.0002299 0          0.00023 0.75         0.0002309 0.75       0.000231 0           0.0002319 0          0.000232 0.75        0.0002329 0.75       0.000233 0           0.0002339 0          0.000234 0.75        0.0002349 0.75       0.000235 0           0.0002359 0          0.000236 0.75        0.0002369 0.75       0.000237 0           0.0002379 0          0.000238 0.75        0.0002389 0.75       0.000239 0           0.0002399 0          0.00024 1.5          0.0002409 1.5        0.000241 0           0.0002419 0          0.000242 0.75        0.0002429 0.75       0.000243 0           0.0002439 0          0.000244 0.75        0.0002449 0.75       0.000245 0           0.0002459 0          0.000246 0.75        0.0002469 0.75       0.000247 0           0.0002479 0          0.000248 0.75        0.0002489 0.75       0.000249 0           0.0002499 0          0.00025 0.75         0.0002509 0.75       0.000251 0           0.0002519 0          0.000252 0.75        0.0002529 0.75       0.000253 0           0.0002539 0          0.000254 0.75        0.0002549 0.75       0.000255 0           0.0002559 0          0.000256 0           0.0002569 0          0.000257 0           0.0002579 0          0.000258 0.1         0.0002589 0.1        0.000259 0           0.0002599 0          0.00026 0.1          0.0002609 0.1        0.000261 0           0.0002619 0          0.000262 0.1         0.0002629 0.1        0.000263 0           0.0002639 0          0.000264 0.1         0.0002649 0.1        0.000265 0           0.0002659 0          0.000266 0.1         0.0002669 0.1        0.000267 0           0.0002679 0          0.000268 0.1         0.0002689 0.1        0.000269 0           0.0002699 0          0.00027 0.1          0.0002709 0.1        0.000271 0           0.0002719 0          0.000272 0           0.0002729 0          0.000273 0           0.0002739 0          0.000274 0.1         0.0002749 0.1        0.000275 0           0.0002759 0          0.000276 0.1         0.0002769 0.1        0.000277 0           0.0002779 0          0.000278 0.1         0.0002789 0.1        0.000279 0           0.0002799 0          0.00028 0.1          0.0002809 0.1        0.000281 0           0.0002819 0          0.000282 0.1         0.0002829 0.1        0.000283 0           0.0002839 0          0.000284 0.1         0.0002849 0.1        0.000285 0           0.0002859 0          0.000286 0.1         0.0002869 0.1        0.000287 0           0.0002879 0          0.000288 0           0.0002889 0          0.000289 0           0.0002899 0          0.00029 0.1          0.0002909 0.1        0.000291 0           0.0002919 0          0.000292 0.1         0.0002929 0.1        0.000293 0           0.0002939 0          0.000294 0.1         0.0002949 0.1        0.000295 0           0.0002959 0          0.000296 0.1         0.0002969 0.1        0.000297 0           0.0002979 0          0.000298 0.1         0.0002989 0.1        0.000299 0           0.0002999 0          0.0003 0.1           0.0003009 0.1        0.000301 0           0.0003019 0          0.000302 0.1         0.0003029 0.1        0.000303 0           0.0003039 0          0.000304 0           0.0003049 0          0.000305 0           0.0003059 0          0.000306 0.1         0.0003069 0.1        0.000307 0           0.0003079 0          0.000308 0.1         0.0003089 0.1        0.000309 0           0.0003099 0          0.00031 0.1          0.0003109 0.1        0.000311 0           0.0003119 0          0.000312 0.1         0.0003129 0.1        0.000313 0           0.0003139 0          0.000314 0.1         0.0003149 0.1        0.000315 0           0.0003159 0          0.000316 0.1         0.0003169 0.1        0.000317 0           0.0003179 0          0.000318 0.1         0.0003189 0.1        0.000319 0           0.0003199 0          0.00032 0            0.0003209 0          0.000321 0           0.0003219 0          0.000322 0.1         0.0003229 0.1        0.000323 0           0.0003239 0          0.000324 0.1         0.0003249 0.1        0.000325 0           0.0003259 0          0.000326 0.1         0.0003269 0.1        0.000327 0           0.0003279 0          0.000328 0.1         0.0003289 0.1        0.000329 0           0.0003299 0          0.00033 0.1          0.0003309 0.1        0.000331 0           0.0003319 0          0.000332 0.1         0.0003329 0.1        0.000333 0           0.0003339 0          0.000334 0.1         0.0003349 0.1        0.000335 0           0.0003359 0          0.000336 0           0.0003369 0          0.000337 0           0.0003379 0          0.000338 0.1         0.0003389 0.1        0.000339 0           0.0003399 0          0.00034 0.1          0.0003409 0.1        0.000341 0           0.0003419 0          0.000342 0.1         0.0003429 0.1        0.000343 0           0.0003439 0          0.000344 0.1         0.0003449 0.1        0.000345 0           0.0003459 0          0.000346 0.1         0.0003469 0.1        0.000347 0           0.0003479 0          0.000348 0.1         0.0003489 0.1        0.000349 0           0.0003499 0          0.00035 0.1          0.0003509 0.1        0.000351 0           0.0003519 0          0.000352 0           0.0003529 0          0.000353 0           0.0003539 0          0.000354 0.1         0.0003549 0.1        0.000355 0           0.0003559 0          0.000356 0.1         0.0003569 0.1        0.000357 0           0.0003579 0          0.000358 0.1         0.0003589 0.1        0.000359 0           0.0003599 0          0.00036 0.1          0.0003609 0.1        0.000361 0           0.0003619 0          0.000362 0.1         0.0003629 0.1        0.000363 0           0.0003639 0          0.000364 0.1         0.0003649 0.1        0.000365 0           0.0003659 0          0.000366 0.1         0.0003669 0.1        0.000367 0           0.0003679 0          0.000368 0           0.0003689 0          0.000369 0           0.0003699 0          0.00037 0.1          0.0003709 0.1        0.000371 0           0.0003719 0          0.000372 0.1         0.0003729 0.1        0.000373 0           0.0003739 0          0.000374 0.1         0.0003749 0.1        0.000375 0           0.0003759 0          0.000376 0.1         0.0003769 0.1        0.000377 0           0.0003779 0          0.000378 0.1         0.0003789 0.1        0.000379 0           0.0003799 0          0.00038 0.1          0.0003809 0.1        0.000381 0           0.0003819 0          0.000382 0.1         0.0003829 0.1        0.000383 0           0.0003839 0          0.000384 0           0.0003849 0          0.000385 0           0.0003859 0          0.000386 0.75        0.0003869 0.75       0.000387 0           0.0003879 0          0.000388 0.75        0.0003889 0.75       0.000389 0           0.0003899 0          0.00039 0.75         0.0003909 0.75       0.000391 0           0.0003919 0          0.000392 0.75        0.0003929 0.75       0.000393 0           0.0003939 0          0.000394 0.75        0.0003949 0.75       0.000395 0           0.0003959 0          0.000396 0.75        0.0003969 0.75       0.000397 0           0.0003979 0          0.000398 0.75        0.0003989 0.75       0.000399 0           0.0003999 0          0.0004 0             0.0004009 0          0.000401 0           0.0004019 0          0.000402 0.75        0.0004029 0.75       0.000403 0           0.0004039 0          0.000404 0.75        0.0004049 0.75       0.000405 0           0.0004059 0          0.000406 0.75        0.0004069 0.75       0.000407 0           0.0004079 0          0.000408 0.75        0.0004089 0.75       0.000409 0           0.0004099 0          0.00041 0.75         0.0004109 0.75       0.000411 0           0.0004119 0          0.000412 0.75        0.0004129 0.75       0.000413 0           0.0004139 0          0.000414 0.75        0.0004149 0.75       0.000415 0           0.0004159 0          0.000416 1.5         0.0004169 1.5        0.000417 0           0.0004179 0          0.000418 0.75        0.0004189 0.75       0.000419 0           0.0004199 0          0.00042 0.75         0.0004209 0.75       0.000421 0           0.0004219 0          0.000422 0.75        0.0004229 0.75       0.000423 0           0.0004239 0          0.000424 0.75        0.0004249 0.75       0.000425 0           0.0004259 0          0.000426 0.75        0.0004269 0.75       0.000427 0           0.0004279 0          0.000428 0.75        0.0004289 0.75       0.000429 0           0.0004299 0          0.00043 0.75         0.0004309 0.75       0.000431 0           0.0004319 0          0.000432 0           0.0004329 0          0.000433 0           0.0004339 0          0.000434 0.75        0.0004349 0.75       0.000435 0           0.0004359 0          0.000436 0.75        0.0004369 0.75       0.000437 0           0.0004379 0          0.000438 0.75        0.0004389 0.75       0.000439 0           0.0004399 0          0.00044 0.75         0.0004409 0.75       0.000441 0           0.0004419 0          0.000442 0.75        0.0004429 0.75       0.000443 0           0.0004439 0          0.000444 0.75        0.0004449 0.75       0.000445 0           0.0004459 0          0.000446 0.75        0.0004469 0.75       0.000447 0           0.0004479 0          0.000448 1.5         0.0004489 1.5        0.000449 0           0.0004499 0          0.00045 0.75         0.0004509 0.75       0.000451 0           0.0004519 0          0.000452 0.75        0.0004529 0.75       0.000453 0           0.0004539 0          0.000454 0.75        0.0004549 0.75       0.000455 0           0.0004559 0          0.000456 0.75        0.0004569 0.75       0.000457 0           0.0004579 0          0.000458 0.75        0.0004589 0.75       0.000459 0           0.0004599 0          0.00046 0.75         0.0004609 0.75       0.000461 0           0.0004619 0          0.000462 0.75        0.0004629 0.75       0.000463 0           0.0004639 0          0.000464 0           0.0004649 0          0.000465 0           0.0004659 0          0.000466 0.75        0.0004669 0.75       0.000467 0           0.0004679 0          0.000468 0.75        0.0004689 0.75       0.000469 0           0.0004699 0          0.00047 0.75         0.0004709 0.75       0.000471 0           0.0004719 0          0.000472 0.75        0.0004729 0.75       0.000473 0           0.0004739 0          0.000474 0.75        0.0004749 0.75       0.000475 0           0.0004759 0          0.000476 0.75        0.0004769 0.75       0.000477 0           0.0004779 0          0.000478 0.75        0.0004789 0.75       0.000479 0           0.0004799 0          0.00048 1.5          0.0004809 1.5        0.000481 0           0.0004819 0          0.000482 0.75        0.0004829 0.75       0.000483 0           0.0004839 0          0.000484 0.75        0.0004849 0.75       0.000485 0           0.0004859 0          0.000486 0.75        0.0004869 0.75       0.000487 0           0.0004879 0          0.000488 0.75        0.0004889 0.75       0.000489 0           0.0004899 0          0.00049 0.75         0.0004909 0.75       0.000491 0           0.0004919 0          0.000492 0.75        0.0004929 0.75       0.000493 0           0.0004939 0          0.000494 0.75        0.0004949 0.75       0.000495 0           0.0004959 0          0.000496 0           0.0004969 0          0.000497 0           0.0004979 0          0.000498 0.75        0.0004989 0.75       0.000499 0           0.0004999 0          0.0005 0.75          0.0005009 0.75       0.000501 0           0.0005019 0          0.000502 0.75        0.0005029 0.75       0.000503 0           0.0005039 0          0.000504 0.75        0.0005049 0.75       0.000505 0           0.0005059 0          0.000506 0.75        0.0005069 0.75       0.000507 0           0.0005079 0          0.000508 0.75        0.0005089 0.75       0.000509 0           0.0005099 0          0.00051 0.75         0.0005109 0.75       0.000511 0           0.0005119 0          0.000512 1.5         0.0005129 1.5        0.000513 0           0.0005139 0          0.000514 0.1         0.0005149 0.1        0.000515 0           0.0005159 0          0.000516 0.1         0.0005169 0.1        0.000517 0           0.0005179 0          0.000518 0.1         0.0005189 0.1        0.000519 0           0.0005199 0          0.00052 0.1          0.0005209 0.1        0.000521 0           0.0005219 0          0.000522 0.1         0.0005229 0.1        0.000523 0           0.0005239 0          0.000524 0.1         0.0005249 0.1        0.000525 0           0.0005259 0          0.000526 0.1         0.0005269 0.1        0.000527 0           0.0005279 0          0.000528 0           0.0005289 0          0.000529 0           0.0005299 0          0.00053 0.1          0.0005309 0.1        0.000531 0           0.0005319 0          0.000532 0.1         0.0005329 0.1        0.000533 0           0.0005339 0          0.000534 0.1         0.0005349 0.1        0.000535 0           0.0005359 0          0.000536 0.1         0.0005369 0.1        0.000537 0           0.0005379 0          0.000538 0.1         0.0005389 0.1        0.000539 0           0.0005399 0          0.00054 0.1          0.0005409 0.1        0.000541 0           0.0005419 0          0.000542 0.1         0.0005429 0.1        0.000543 0           0.0005439 0          0.000544 0           0.0005449 0          0.000545 0           0.0005459 0          0.000546 0.1         0.0005469 0.1        0.000547 0           0.0005479 0          0.000548 0.1         0.0005489 0.1        0.000549 0           0.0005499 0          0.00055 0.1          0.0005509 0.1        0.000551 0           0.0005519 0          0.000552 0.1         0.0005529 0.1        0.000553 0           0.0005539 0          0.000554 0.1         0.0005549 0.1        0.000555 0           0.0005559 0          0.000556 0.1         0.0005569 0.1        0.000557 0           0.0005579 0          0.000558 0.1         0.0005589 0.1        0.000559 0           0.0005599 0          0.00056 0            0.0005609 0          0.000561 0           0.0005619 0          0.000562 0.1         0.0005629 0.1        0.000563 0           0.0005639 0          0.000564 0.1         0.0005649 0.1        0.000565 0           0.0005659 0          0.000566 0.1         0.0005669 0.1        0.000567 0           0.0005679 0          0.000568 0.1         0.0005689 0.1        0.000569 0           0.0005699 0          0.00057 0.1          0.0005709 0.1        0.000571 0           0.0005719 0          0.000572 0.1         0.0005729 0.1        0.000573 0           0.0005739 0          0.000574 0.1         0.0005749 0.1        0.000575 0           0.0005759 0          0.000576 0           0.0005769 0          0.000577 0           0.0005779 0          0.000578 0.1         0.0005789 0.1        0.000579 0           0.0005799 0          0.00058 0.1          0.0005809 0.1        0.000581 0           0.0005819 0          0.000582 0.1         0.0005829 0.1        0.000583 0           0.0005839 0          0.000584 0.1         0.0005849 0.1        0.000585 0           0.0005859 0          0.000586 0.1         0.0005869 0.1        0.000587 0           0.0005879 0          0.000588 0.1         0.0005889 0.1        0.000589 0           0.0005899 0          0.00059 0.1          0.0005909 0.1        0.000591 0           0.0005919 0          0.000592 0           0.0005929 0          0.000593 0           0.0005939 0          0.000594 0.1         0.0005949 0.1        0.000595 0           0.0005959 0          0.000596 0.1         0.0005969 0.1        0.000597 0           0.0005979 0          0.000598 0.1         0.0005989 0.1        0.000599 0           0.0005999 0          0.0006 0.1           0.0006009 0.1        0.000601 0           0.0006019 0          0.000602 0.1         0.0006029 0.1        0.000603 0           0.0006039 0          0.000604 0.1         0.0006049 0.1        0.000605 0           0.0006059 0          0.000606 0.1         0.0006069 0.1        0.000607 0           0.0006079 0          0.000608 0           0.0006089 0          0.000609 0           0.0006099 0          0.00061 0.1          0.0006109 0.1        0.000611 0           0.0006119 0          0.000612 0.1         0.0006129 0.1        0.000613 0           0.0006139 0          0.000614 0.1         0.0006149 0.1        0.000615 0           0.0006159 0          0.000616 0.1         0.0006169 0.1        0.000617 0           0.0006179 0          0.000618 0.1         0.0006189 0.1        0.000619 0           0.0006199 0          0.00062 0.1          0.0006209 0.1        0.000621 0           0.0006219 0          0.000622 0.1         0.0006229 0.1        0.000623 0           0.0006239 0          0.000624 0           0.0006249 0          0.000625 0           0.0006259 0          0.000626 0.1         0.0006269 0.1        0.000627 0           0.0006279 0          0.000628 0.1         0.0006289 0.1        0.000629 0           0.0006299 0          0.00063 0.1          0.0006309 0.1        0.000631 0           0.0006319 0          0.000632 0.1         0.0006329 0.1        0.000633 0           0.0006339 0          0.000634 0.1         0.0006349 0.1        0.000635 0           0.0006359 0          0.000636 0.1         0.0006369 0.1        0.000637 0           0.0006379 0          0.000638 0.1         0.0006389 0.1        0.000639 0           0.0006399 0          0.00064 0            0.0006409 0          0.000641 0           0.0006419 0         )


** Transient analysis **
.tran 1e-07 0.000642

.end